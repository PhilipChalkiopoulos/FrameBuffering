��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�KW�UHս����fP��nIw@��Fn�~�}��w�{���ڽR������_^�p��1��q�ڪ,�S鄄(I��jx}I�����y�"˜idW\��9� ����l/8�g�UB�Ə�7��s���#���&��4�Ũ�/�85FLHE�t�)"!�}�F����L�AfY��I��I�I�(�I"u����~�t����_�ʶ`�R漖��-twz�S0����R�	ōU�ّ@߃g��Ϊ���|4±��P�Ak�gvQÅP1��p����4����=�_��j�l8�5�\��6xc�����z"�����|���!톼[����g>o���;��W�yM���M-.�E��4��r��ve<j9x�hL_�
��Y��O��R1R�����~���׀���u�ަ��b�,$���}�C6� ����S�w&�A��h�3��,9����KYo�[�b�E��$�`��t*��>6�� �ć~�����k��Pe�����	�M�K�����~�*�ʆ-P�ss�;��>8�[O��Ǣ���Z���+��-DY�����r�;XdR�$�dQ����UI2U�}>@7S�6��Ăm�Oև�,���3B'����1o
�[~��MG��+8�K�]�ߔ>j1+�O��->I�k�y�u$�+S,,�M�kq�j������W#T�'�I͏��A����<�����t� �K#?�zz�{���@���1pJ��}���jdza�
���R	�]*n_�JT3��z@r��W��le�z�e^��V,�v=��$�-���zɧj�0C`z��[[b!{�E�$�:���<�����IB+*������ŭf�<Iݾ����������$dE�M�wO�}ĿXťq隬�z�0l�e��n�����B.�&�j�[0E�	IT8�����n%�ˎ�	-�O�"��ގԚ��z� şy��m+���P��n}���C�\KM�DoK�W��'~F)85m-.�_83]e�eA�'��Q��i�vL�Ƈ;���P�#�3簿+�I2���!���p�u�N��$p;�.�f�5QB5XMs�(�K.�ن�%��f]�ia�f�M���d>]a�q ���l���\��������l��Ƿ��p�b|}����1sxJ˞���$��������p�i}��� |���^H�p/]@c��T�W�0���:5I89�jū���� <^���g���qB��w�qE���6ױ~��T$�~=��K��̓��KF)�XIg�x
���f�p�r�;B��(�;�Ę�$m ��_�&<0�G�ݦ#�X?�W��L�t��{���lJ��+I0�
�m(�e�v耪]���;�\���1�˄��WF3��+8�u����U�=�[/�o]��$d�x�T���4c�Q�,0���u������l���ɫU���'J����;��: �ۇ�O�����I�#_�T�|+˳�L�n}���eX����>�5n�O��)��'�^�
�������4d�.�(��"보��#f&�X�2�ȗ+�Y0���)�Z��ق?̅�h�Ӊ�|�(���A��,�N�2I��lմo
���o�f�dC�Z��/m��!���?5���'��0"�ʄ����󱦎1���Zʶ�J�#�=�3��J�4�Q��>��n���J�X��1�˕��i$�9k];�7�[��C�WE�nbD+MX�����^���t�9>y��g�� ˯��">�f�
ֽ�b->��K@��Y�U�����3-�=I�*���:�V�O;tJ��.�i;Z�%HrlnXf�!���,�%OA#z#�d4O�"G������,�g+�Z`�#��"��:�a+R�=�>�jc����CmP��#1�y��g�x�ς�o�w�I��C4J�u� ܏&�!h���m���g>�,��1�`�!pK���7!��{�o�E��g,٫,�g�ݏ�b*v�\9x�ݽ>��W��U%��v���^�ֺdd���X����١Q�Rǁƃ=��ߋ����6
��A�WaPU-����О��{ _Y>�5�p�����ua�2Vr:���������j�Y=���[�Q��e+\�D�\�SS\��x�p�e*+���C!��~̇b�?��yx7K4ɦR��N#aē��p��N�25�8�o���3�zvW��c�"�x�MEq˶4��U��0gNۀ'�u['���S���H$�1kmͺL�Z�ƛ��5G�Ã�އ5�'�$�6;��5�]��������R�͝[�{����!��0���?j�xc`�}�kmH�M���ޱ���S� �uxF?���(���� �=��V^p�]8����2���'��)��3u�Ǹ]�Zz킐W!��ip36��G�D�����VvBw�r����~�5�S�\�j��`ZR�e7Z_�=1� p��B�h>��d�-�=Z��tS��D�L���Jމ6>Q����������?\��l/y��y<$a�ɳ!��P,߈� ��C��."��I����s�e��Ϙ�C�2�Q���ۈ洿�$,Å�Yq°rh?F߿�%|���D }��k��1�6"zZ̢]:�pRخ�]�h#
��{���d��o�A��ֳ*l����|��dQT�l0�I�0��t���HcC��P��Gp���|������Q��brϝ���M��������Y�ܯ�vY���k�������#�����Z�6ɉ�/wO�;�����Q�Zr�1q����R]��ajj��H����
0%<��9��K�Qy2�6�
+��1Ui�!��J�C�"ѮO�� �����0,�y�ţ���ٳU�h����z5I� �q)�z@�����2
��rb�zJ�4&/u�c�z��}f;!"!"��)4p����N|�AX���Ԋᾳ4O�0K�M�]�2P���^�j�6��l�гi�����7�!�d��,VK�S+p��~��������b:Y��J�
�+�@_� ��yIa�BN�쏺���~��:Nq��B�-P|�˥;�/P3��j��|�.�����#$+Y��jꏖ3�Ֆ��-N�#?��������~lK)�,H�iD ��S%t��Q��OPL����? j�G�%cm#IRR���S���9����Y�JaƲQ0�������V��q�����<��O��E7k���\�������4�����%�V��<�h=hh�D)}w׈� +�$\:�Ms3�x�m�6�f<��p��62�Wd4���^�i��f)K0�q'c�~�PR�f
�Dx���F�> :#nunB��Z���ta�k#Ƃ1]�����-J{+<k8��&�<�����������ӆ�������ͨ�l����]~�R��f�޶���K�d����둸m07|D�2`��9���q�w����p���pXR��_���)ݬڄQ�`m�r��0��k��A�9��J�z^ҽ�o��#=�R�ߵ�T0�S�;u���Ʋ����cUw����Ѓ������/�k4	ְ�@R1k	�+3Pd3T}�lUA��t�`BS7�gV6�.�LH���%�t,�7��󺼕'Iǥ�F��� S�$��{�=&�[�̦D��r,�&!��S��A���Mkw����TfuRl��}�҂���j���<��^^UeF %�m�YSJ��#:p�gx �U�2F�����H�\oV��LK��4r�&s5�ar�DE�Q��Z��@O^�\%�����z50��С���!��<_��<y���%�Xw��ض�^����	u1&_k���*�D4؋\�a޼�u۟�%�@�!V�u��-�j�HFM�wg�tw�V�5UD4#�f>�H��RB�
7,CZ|<,0��;���c����.�7cӇk�("�w ��ӥ�LI��h���ƌP���Y�&�|���g���x�0�%~^z
��L�� �Y��o��;~����5]�O�s��.�ӆ�vnԀzN��KGY� ����#�d	Yp߯��c�13V.֡8bkTt����$ص��<�n��vVR����{R�)�oP^b�1{�8��eu,�
.ga�a#�Q�v�̕$�+m���ys_��
�ʊIm ��6�՚��+!������l6�n���Q��2{ݎY�3נ?����\ ��o1��g�2ޥp��en50�Wڕ�����Y�Q�MG�7���rD��H��D��(:ѭ�P.}���(	a��D�}9U�/�
P{��+�W���;*�$:�J�/&2:�ic�.���лp�cd�_!s[��+�[�a¤���^�DaoTQ��T@�R��j��_3A9�É�X�v����͛�(��wE5�Y&*#�=Eiv��i�p��E͉cM��h��7�)B��q�j��7��{�k��C����>�o��ϓ[���G@gm�Y���\z�:����1.l�xxӺ�.�|ʸȍR��Ӡȕ������<�vD�q�z��:�����c�T#d���9��E��� ��,1��þ�G-<ᯞ�����g��A|�0w#b��2���a~ĚH���z�bX��|=�L��*F���5�o�[q�P�S�����԰3����@JR�v�c&�t��08�B�)�xD��^�4k�����c�j;��Զշ�)0�C��?K��p�+T�6áo��15�Fl�0_�L(
srlZ�@>xK���]I�X�)07���\���8$:S��R��S��!"<#�G�Mfo
�|#6����:#4�?Ǉs���D�ؿ��Sj�*����ÅBS])�xӥ��;3�r';�������|}gfĞ	�ʞ�����ʔ#���oI܃)q�4����g\���_s��f-��)�|-?��# �f��v��%i���H�,ɧG���4Hڐ�ks���4��j!�0s>�����@D�R!�b�>��{r�A�V[��C���"
��QT�gbݔ�+UZGm�R�$�T�"�Ǟ2Tw��1[���<|�HH(�oV˭����a���xje	t�Kt_���e�/��6�e��Ʋ�>@)��9pܐT�N1�fl�zG+q��Z��W>�\���l��;3]g���t˷/LpA�گ<"/����l���OM�֢v�P���Ś����e��Z
���w̲�J�5*I�_K<��>��$��#����=��d�dT]�fS�=Ъq��E}�'�����K�)B,2U�1�K�ԛ>�:���3v���e[����<��Xn>�[��,��4�>���|��9��M�ɠb�#�fDr�� ��G������F���!�%�x��^2�P$E��_��&�(3q�|T����X{��!�g1 ��'�|�!�w ����+���|��1�2i�q��kU��+�!7�U�C��%
&8W_u�' �mj�>�%'�-"����?����� �3$��kv���Q&��S��0c��}r�<0����������O�Z��+[b#������Բ|����кK~F��Jm���z$�U� rb*S��0�J�@Y�������Z�<���	 8�߯Su�
7���ge���``��6��<U4J�%�a�	�T�a������N$��߅+F��k��j5=��n�S�(Xb����Ћ��r�����~ծ���%�����|��	�:���������;��d�{ӡ�Ӻ]d�؄,W��Q��M�f`%��ᔽ@ɀ�H�K���#��:�+�:��+aꮇ@B�Ɠec@�����讆���Uxɰ�W�����F����s8D����F��ݞdJ�����C�����g�[�{.)��əđqΘ�{/e��#<����U0m�mv�{d�N���m���u�1�+u	ɘ%w�A�p݋4h~o�v�%ސ[{�Rn'e_$E1�L0'���L���-�W[��5O����3W�W(�.b���ޫq�Y~��wnA����0~�Xü������QP����{A�Eܾ]
�cf��eKB��j@zh*� � hD�o���@Er�a��^�ZO%�=����}Q��w���KDұ�JA�?A��\5�)劣��k�"��ݹ�A\O��Y��o���NC�v�x�[�,g�x��)9����ݧ�`.�
ˀΩ�Ȯ��1Hu��h�Y�z�hl��N���i-TX�@?* � ���G�?�
��*v
�j���Cߕ`Ń��^�`�����G�|�lKjM�I�3�]�!�8=��T��s�EaGe%���R����j,��e��4-���	�aPF!����{
�6�Y86���K��6��rĵ?��}s��h��Yە[��6�8���梵.���E^t'�.��r��z}������|��*��6Sʨg�����$���P�ʩ(�}��mGf6� X.�'�������;� ?䕸�<M��艿d��a�����&�H���=,��?�w�?�~�3�j���O�}�sk!!�h�Z\��C�`�ǆ�#��I ���M�,����D�����f�d�#����[����x6Grw	�����?P��,�k|�J�{|_�9?,�
&����B7��Q�����>��r��e-���8�i�ޛEؓq&����[HT�b�;�@�Y��H���A�Ҵq���ϝ�Ԍ.��Ȑο�"�;��%�[ι�(�u[�O�A����)_ �h���O���[��6b�m������
L.��+��O���`�ެt����ܼ����.%�ɼp^��WD߱��L/`��5:]��e�fEq�0�ͯn8AB�\��p�E����}$?�'�tgS�J�7�@	�qe�����\o-�e�3![�f���܋�6��m6%��]���4� �L�t�4��T�0A����ܮ�ök�p�|�p$���=UT�2�������b�_з Vq��i@q��,�ll�C��Ho�����Û�L�Ӓٲ��͌�!�[E�GeƆ�ً,)(�#�������Y�d��Rjb,$:߿�J��G����nm�u��E��!�/��s�4'����r�]��q]����
�H��y�$�[ڽ�.KP�)3���a�������	��Lg8�t}�Z'g4���Ж(z7^k��+�6����T���帓�c�K�s�����]b۰!Bi�ۦ�{sp�/ZeJp3��m@�o�f��%�����/�Q���5��^g|Vrʑ�P��=��!2���䡘�L�7gtMI��M9z-��Nff�F��MغL�18�P
��*}�Fmѐr\�x�*�`zR3~VO85e����5�D�p.9&�̽�)�p�=���q�K��A]�,^,�!eoӊg�U�z`�\*M����^���*���M
���0iQ����p��f}�V;g-q�{�I"��� Q&��Q"x2�#�v��&+�u�[xC ���俎B�Ujl\1�cyO/CҰ�^�;
O�Q��Ͽ7��hh*�t���Rk�FQ�5���;�QX�!�����G�Α��3j~�}�uq&��2��!e��^2B�M��'�t�n�b�:��̑�v *B��%E�t��v��R���N.h0�F凜:� !� ��N��є���z��<��k/7�	T��az��먖�>��J q���4� �c"e�`�,�}ާ�Z��hi+�,k��U�Ȑ9����P�=�_�7T7�U#ȵ�y�Qߖ�S��w���?�X)���9~�fwb��+"~'�.����������A8�L.s|	w,B�9WQ�" ����NOk�k�;Q>���X����(�.�,��S1Q{��y����F\dc�Y>���:LLZ^��
��y���K*�bg�$�p/M=���ߩK��R���M�'Gp�0�y�U/Idb�e�by��y���W?�K��+׭#���=�I�a�14`�QNz�M:��h��f��t0�����q�D/)�A���6��py(����9����hW�.�br�� �"��|M���I�D���iD��:�+��,D��-]n�d�+������Cv���95w߃�G�\��_"z��"^��9ٜ�<���<�%�v,D��|a�|jLer�YP`�- ��#�/X8/k_ȥ};���;����~�Ғ�[�uvu�;X]@�|�.qK�وbf�b�7���m�?C"�!�K��ߔ�.K���.�5o�I'�u>:e/�;�f���ރ5&�^���d���	,�prV�;�-�L{o�Q�ɧ#?��~[>A���^Vfdz��B黰�)}g�쳖P�{��)���R��U��4���qj6�ȓ$���-��kӅҠ�v6꾅pC��[������('&fx.$�}�P�${G�&�QNn�%
xc�>���T��WS}��^q�s�Q��m���A��f��b���s���B��bKX��掼9n����FlU��с�O�$�k�?`M��c���g���)����u��h�X���Rk	"��r�)l2��Q��x}D�ŧ�JU�֫C��>�҂��g���2G!d�bEn���i�J�����y�=D�+�@��G�v���A����I������`K��x�;͑><e ���K �6C)⊢�5�f#^uZD�6+?	־�Dڏv�������!�Āc�0��H|��D �L���3H� c�oέW蝅���1��6	�JH�Rթ�vO�,�I��Zm]�;���`2ݍ�Sj�����z9�zL	9��D%��3a5|\8�Ѵ��~�t�E��'��~x
9's�E���߉T�b�}���w&Zq���LZ�Ht�������=��CaQ}x#L�3Wr��J��a��:���� �Y�Rh[�{�s�S��g�!��=<#E���w0��U@Hr�>I��:�l�:ˉ�9�o�c����0���8�ט.��T[� x){����Qn��V�O�GAN+ͽ�c��)T4����~
�˥l&�g�~�k)�	�#���.R..s��1H�������i��oE��	�)��#B�+����R����p�T�9$]��<�h�B�S�F�Gla��x<�d��c,cُ��O��;��UE1�o�"�'�ӵR�l��!�{v���d*.���UH4P�V
������jM̳��N�p,C������(�:j�=��}6���x����ճ������ǐ�y0n^Ll�"ʿҴ����-��@���Qcrz�x���������P�t�Bj6�9���r�}x�(U��4����Q��:��nڧ���/�!ͺ.c?-��/��}O& ��M=%�ɓ���mx` k�v[�S�.��<ŏ�1_�vB �g��
Q�N&����	�.U���9�?�_�z?������-�#N�3ME��o`ܗ�Me�G�}]��5�x�^2�-�b$
`$$i�7+�?˥hձ��NG�R�H�VL� 0���5�.�d�:��%w�C�E�}Z�W+fI+��I�����/�U��w;�H�����ĸk��+^�����5ȇ�?���K~�3WU��[%I�7@�6�-��?��&�^;*K�b��;G����� �08d��gs�E��7����2�1�N����}E�洺Z�*�� �د]��3z���������H��6Ѳ��{��ִ◅_ԯاf��R eۅ�������$��/ۥs-���l�1�+��(x�9�'n��Rz��	��3Z������1�Aw�PG�t�v�>t���}�m�u���N�y'N�`�?l[���;�G�6�͸¿]��m�乓����I�/g2.{bl�t�C���2��񻢱5C�����H�w=����TV��Q�~C[oxP	 ��C�e��67��A>�6`��6�Y)���� �O�U\�psFf��d>؈,,� ����vf�K	4g<Q��9Z�3$����I�x��/�h�	g�5"��Pi� ��tlټ���5>'�#X^�K������Q�r+ě�]�e\ZEH0�����XȰ��m١�@��rY{��f�������-�<�Ni�p�۠^ݼL�M4��XE�h���xn��^��8
����?p<<[r����Oj��j�<�����Н��;��=���u9��Ca:�Z���>1����1��e�`��}�D�߸�"F�q�t\�O�`�Hd?}e:�/mol������M:����*,�(נ��U'�e�����*ٓ���ii_��'v�Rxms��������~ ���]�ڎ�د��4h�<�5$`���N�
�6�Vvq9T�����ưp���Dm%=�r�V+��l�AN�����-w̟�V%��2�ٕ̦;�/�@�t�X�B~���������	{r�0Wk.�Z�g�[���{�Z��xz<N�m���l:��E���΀������;(�htUҁ�M j:^����:�8iK�^%;��������mR�Jj�x� 8����
���;&�j�Y�q=�2pԲ��_"@a��d���h�ւf;�Y^�up)G4p������uG�y$�D�8=u��u�L�OY�S�J��k��(����(0����B��o��,d���᧵1*k�;]d]au�i� uąƶ��u�i�=_�Q��wa���[��P��cx2�A��?\mS�D������#<s ��[��Pe�LSN��X�8�7�����d���ˣ�_T<���b=�߉t�^��N�瞻g�{<џ>�r��PY{����'�����S,TM�paW��H�w�����S ������e$U^���vnxj4P���IS8��L5�_ny�{/��QcJF�OV	1����jS["7�k��rh��`w
�.��� -�����_�M�\�:�V��ID��(՟�NKAI��6M̨��yO��	\q0��x�H7���'��)C̜�#1�[ŕ�6�,#�k �6��W��h{�������~��u�Sja�Pq��t�n�Z�]a�q�m�gg�t#P�u-��"��qA�\��U=Rdm�5v߆�Z���HP�uг*E�EY�u[B7}����x��#�iӝ��]��q����,_ ��R�,B	�JkW�d��A���L��u8����D�o���┚J��mT�%�DV��{F�j�}����[e��t2�M�4�ʬ@���ݜ�!5�����u:�jQ��"r�IId`[�%rq��g����dd;l|���W��O_~�0ɷ�N����^*�ؓ�L���A�ǁ٠pţɶ����R���EC�9|�9�x$���z���RB� *C��W��e�B&a:;t��e Cu�X�8mR��F�mn~*��Î+�� @=8����P���c�"�&��E/���q�j�\#�[ښ�Tvs�޿�+�ʍ�*��9f�g���髿i��~�=���Ʀ�roB���kM�:��AC�Í�+ �� �t���kuOj�)Sm�m�"���vt��,zڝ�A�;K,�epŪٰ9��S� uc�=�����3�4 �=�ӑ1h���Y��4n2Aa{�1���f�p��K�;Sq&���~#�y`[R6�[ԝ�An�F��X���N�c�l3*��]��U?�P�e`Rx�_GS�ud�d�1P�f�`�шs�0̄o@׫�m���a�A��!�޸ef�R���1��3�;�XW�"p��Mw�h�U�rJ4�Ns�ڳa�Iuo�R�p��'J�͍�����2���Ag�c��TLwݨ�cL̠���ܖ8� �XҴ��TVD��ߺ�s�K��l��h ��ޡt�c�fn���{�ߏ�:}���'L��u%4_��@�Vn#�P{뚽�SL�[����g��ضLG}�x����
��j�7~��@J�ا%~q�	1���1+1����}�G	B�R�J�DAd�,S(?m�bq�x &;�]
K�E����Kѵ�ẻ{ �C�
_�Z5]Ak�<g���t��+`LM���4�s��~rW+�� 9�%���{���L��2�KF�` �>c�1$�8�Wq3z�j�������0�phz�Ƹi ����ђ���V�������<����rBb�u,Lj+H�X�I��m�e�� ����b�j� .=�$���`^ي�Lb	��Mn�t������a�9�n}�U��S(��c���Ji&.�^�_$�6���8���ޡ�%|�Q����s6���A7~�e���I��+�"3(��L[�։B�3�{<�7	�a�O��s���bP��g�@��n�		\�T��$����9%l��ߞ�1�!l�Ǉ��%h@�"2����
-� '�h�F�W�V�V���3lZT�ӟ��57�J���4�SO�$��@y���+r9��F^��L�2}������Z��ц��YzL|"�j�q���> X��V+���(@�)wG�b�'�����Gϼd��Bީ���^f$��;��߽G� ��KwOh���&�x�f���9H����QlZ�d�䡃�ȭ���)?<ɗc��:)l���:7&�����'�?.#�k��_Rd��N'�c�B���J���n�j���YU���}�27��2���8�=�i�*����S�De�"Gط; ����ѹǅ�����N����(\Ut�(�� �b���j�CR\��hFX�80���������F�/E+��_�n��"1W�Rb�N$*�*��G�Ky�s�<�A���Y!�WP���n��+j±�kj�;��-�:#V_��A)�q`L Ʀ�X�d�p���cE�6�Ǵ��������%�i����u�Scv�#���C27�U��S`�g.�\HO��q�}�d1���`>)�$�mdv�>8��0"I�%7�E}�M5�v�U��Ac��ֽ8��w���&i�
�,�/#��%�12q�#h%L�eeq�H�p��L�&�ɺ��Eŕ�o�3Ɣ�/Ȯ��Ƅx�u�I�~�+9�$y���XHrȸ��2F#S���{��� ��b$2�pT"}�h��m9j]���PN���f�j���gPr��˫\���E���h�����=X3�j����l��O�i$����{.�X ��_�VR�.7~l\�Xb�%x�'��h9�o�q���yIٷ �sF�NC��tq8X~j���Uz��n
�
�����t�$1飿4����՛���mY�أ�J� O[�A:K����o�S�{D����!a�9z6cUC�Zy�#��4z����j��[�Z�Sl���J��2����[pi���9pF��=��U�}d��Dv�M/qLϢ%n�jР-|6Ͼ`&O �b���6���h�yt�[�L�Fo��/��y� �֓�v���3�Y��
��2�(u�Q�y��jI��Y�x(K���M�?�H�k�yJsXN������+g�ә㬦�O��8z����`
��������乙t�w�[bج���u�p��ඎ��g�[�Ah�T���g�Κ-�2��#g��H�#�pBwbAD����Y����X�C��kG�[D��r�pPv��$l�w�fP)�0��7��8�
r���)�����ƸI�H��D�Y�9w����r^�P�aҽ�x�an�Y8�}����w:j�J������fރ/Lܠ�w�P����a�1.\�>���G/���0bĞ��e���d��Z||ӥa�麟-��8N�-��_�N�t��y�*�����y�b�{`W��\��S_C66pĎm�G�����&��8�Lr�6�k�I��ʽ��i�% ���Z�M��Ƿ,���rKݕ͌3�vu��Q�^%$"�������,#�����u��6:�钔aY}x�~�0���%蝕�*)`�+�HژP�����ꧼ��L�g|6���?%+w�
���+t�����A"�m~k���*�ְ\Ĺ�O5�<*�*��O�Y{^��x3���.�+�FǞ8e�y̠����^��5�������:�^���&�	n9i`'m��.|�rӴ�����b=y��v��x��>?�ߵ�����Bj�>JZ��xF�����{/�[�"cZ� �NU��p�@�\T��������[,�?�u�n���A��CK-�h�s|��D�ّz哜��<K-������e�^��9����!ᜳ1�����I�!:��r�i��{N;Ž�uh�Kt�5��,e��Ix�Oņi|�
���4��פ$�n��>ﭲ�2�qρ�aJ̶��	�˻i+ľ��u�Aiy�	7�-���:<��{��z4q����= �/�Q��4@f�Sf����X��u̬[6p��Nm���*��$�I)���9�ېꬮ�9�|96���jvv��+_���J�c�j�TZOY�����Y@ Ecz�eT�W�kk,�� aa7���e����h����$�Ac"j�4��]q'Sp���Vf���s6x��9���.��0]�8�*n.�p�E��Z5�X���������M=�[ϸ-��D�U��b���4���r��H��j�# ��'.�bj��x�d�e��<�n�_�$#i�� 1+�j
<���U�w,ʅI�.% \N��=�&?ͲϺ�A�ݪ
����(�r,k{R�����?��̹ B���#�z�� ���A��W�d���d�{z�/"]�3��"�iQ�����k�%y]����/�+��<�v`�j��V8 �ϱ$����u������qe� 6�t���2.W�����>�T�P�X��+3����/Bt�֒��j��j����vm+�G�#�]�d�ȟ3?Vj�0Qf�̙bх�d����'|m�aݒ�»v�(���n������]�@�f���y���uPS����r梿�l �������0���yL��	���V��(����gNv1�!l� J��*�[F0����2�_������d>b��D�^e������������#�����Cը��:$*�6Ҫ�},Ƅ)4YIi\��p��\gL���BI������5��tʬ��4�<}�R�sl%'
zÉ3�W-�T��ǝ:Z���a?��!Fd|4�Jt��[e��&Lc������d���E�p��	3kj�7A��"��&M�k����-ҥ�	^/�ą�b���2�G*vA^<np/ �B��%�(�n�i��/-�
(�a��X��ϥ����|��\��+߃.�Ц2�:�lp��u�r���K�����}��,�R���9wW���@�@x�H�%&!҃7x�@�݆ߪk<ƚ�1�85��N��}�@bõm4�p� }8�?	�xڴ��C�e\�9�l�q/��@�'� �f��;��.�א�w
�J��!�pԸ��į�*H��Aׄ�,��뇿�r�|�U��c�G[�_���#Q��5�AAk���vB�X+HM�c�O.v��3p�o}W��] � x��H��Bm����^XRݮ䇹r����ϸ�� �\�Y�ɥC�.aW�A� [�ƙ��q{�?��g#|k��7�_ҹ�n@��1�7�:�43Tx�v��dhz��YMv�4<rx%�5}�*����0�S��X'�E�-�M�&O�,\�g�g��T���L�������W��d0/�b)�@b5� vj�
�+.v/r���e����tg� �o��	�#�Kvvɡ���A@��:�j���$�y�@����!��t���v�>ĒX�д)F'A��;b����e��������%,��348�����ְ�aGX3W�g��63 �b'�)�:ա3��#�S!��H����ۤ^H%g�A@p ��켈����?s���=Z�%i�@�J���T'��r9e��t�Yq�n$�e�^�Fv!z^�b���m�^?c��q�Q�=��V����C;�����"�o<fpB��Br%˂���(����W���\�`�����M�k��6�5X�LBә�ͩ�؁
�J8`8��ԡCj�xL�:���m��*w���Pш=��_>P���{�nop�/�1�X��v5���)���g(n���̝�V�pH;!�����B�&��8>;�ʣ&���Ug��R�E��͉�@��>H=?�y=ff^"�E@fe��y2�A�����V�~,�Fey�(�w�ˍ�.�J'?۰&�m/����i���8_�;1��$3YV�a4����@:]�+�9�R�;����}B0���{�:0���|��� }�e� _��7ҷ'�|�g�:Xe-GH� �2x�"�ޖ�
������p�w�ա��=����H���S�����4�NX3���""����9�9`�F»�CPK�l<�����T`���h\@�ҁ�2�V�l�<<��9BBB߫��J���\��Az���*$"�εs��F�2_A��#u����3��!-��i�v�Q,��*>�ib���]oB��&A�Q�Q�C��1@����.�\�U��?$���	H�U4]��A�37ɘ~2x��W[�s�ͧ�9��96F9��OS��ѯy��=7+��`�dR�P��Q,����)�Ŷ@�xg
PA���đ��w�wl�_Rz ��7J��-X�mq���aLe��t�ρ⬊K	������I���e��^��������`�k�E��;�:�u� ="���M�P�)��O�V�9?nK�
�ZYCw ���'��}{��c�4�9�����9�-�^4�����l�/L�Evמ�.A�l���~�zR�<��y<�L��&�l����c�A�I��I&S�@���K2C�|�d�~yZ��Y;w[O�@�̀�u���/TC�	̗�і�'^�x�����9��:��T��.�h��g��>�޾3�;���W<�VU����`sh~[cX�*�������e(�- ��:8D�F|7:OgeŹ�EﯣQ.�YNY4���L	z�9�����+�m�2+o_�xh�s�j�4��G���]CG+2U�������{�)��5���/ڇ3*qkԨ̵:�w�@ˌ�9Te���e�bha�ډyTE�0�2�G�� ��f#��xz@��)OW����p�r�t#��v%��K�Pz���.�C�x>�L0�0�.�p|_�֥�����`03�Q؝�N�ݷ�P ����V����qĠ�P�-�������&@�������fc��36YLX(���e�`���꒨�4kZr��0F�aθ����1BQ��]��,:�}�k+U!�ƠPd�妉
h�F�cc� ��m}�P� M,� H3)��?�G) u(o�}X�-���\x�LU�O��P����,��Nx�m�X��,ɰzu���x���0xӽ����!R��m��}5�YU�97e$�T?q�(Kr"���2�v�"�_�ߥS��5Wy:t�n�x��kd�Ia�%A8$E���Mױ����H��Ƅ����D#<��Y�H�i�T녟��cD�|�0�d�7|��������q�Zw�m<�j��ڹ�$܍�u���؍�c�9E}�����[�2xrv8�ʢ9RC�V%���?)�uo0��ǕW���QP���9튳�;����G�\�'ũ{N��`-����;�
y��{-f��LF'$H�"֜����(;�.Y�b؁��Xv�:��P���g:?ͽ�hfft���'�!P���-/2K�c��ݪ78!����9R�M?�2"��N�'
�B��;{&���FWu� �v��SK!M�Q��R��W^G��o�fh�H'��GĆg5$�#��w��N
��g��sq��P��wFá�`��(=�Z2�)��]�?�
ˁf��z�����uD��&��W�`��l0zyο:�*F�6h�30�t���P��E �ߚ�F6���qR{�$����[�?k�ܨ��'���Ph���F�{2N��$ޭ��C���Wy�0n��k��*��d��pGr͛kTz�`\Bf���:��E��� %|	�yP�7/�7��!�A��U��H]��p�����ҍE^k�=��3�N�E�i-�IA��r�#�KIe<0f��}�����u�xMs��j�!�b�ʁ����7棾�E�wZ�u"����>�ZW���_��hW)�=w��?nV(�������	�;W7�c"&\�!7A�F�U�?;�Ox&T*��)8���,[dkf}�\cjO�C�k�7�7a��4Iu���k=-���]W��cC�k@x������XW����n�$�#� e<c�v�<�a�ȷ���f=�~�����D*"���;n��/��:WZ���%��pcJ���nІ��Q�z�HO���a��)�ڙ���2���g�;��h��ӕ)Gm� ��gB���Qny��SN���AZ���u�ե># ���E�۩ѝ�9G�/���[jA��M0� IY�m���3�Ӥ�S%���������)�%,b�Zbʟ��8��[o�5�� �� O�[�*�y�A�RÊ�'�(�:d�[DX}9����t��������~d\�=gw�:A:%�j�-���Oi��9��
���&D'b�hN��e�a���������j�ȒQ���0���"�aZ�DW��H�y��܍��9��S8�=�<��X��B�ǥ�
�:�$����8��6J��B��1�j�M�>���mc�(1�X� �~ր)^�h�\���GktB�&��7ז�A��9��ˎTl���mW�o>�"K8�D��yR/����IH���¸���(g�2/ݙqBS%���Xu����E�
�ay�[�u6-x��4H<��V��Z�~�|�\��@~�s��m��?k7[����ؿ�N8�l�uH�����j�.�%��E��o�"�='�t�����U9���M���}�W�|�˜���
V 9���u�6��&�:WqH��2��K6�T�~:i�k�U�l�}E��0�b�>6Sϣ18�	�)�(Y*���U�7���*�K1����m�>ۼoS%���y��?����s��`��q�K��YX�in��Cu���� E<��)��jpe���M�����L��9���A�.��;>-,�#�S���_�Tpj��j��Ǩ�{��[�����Z�![�����u�z�N<�R��}C0���SB�R~B=���IcK��}Q���5����u!N	۸AO�b�i��%i�ݿ[P~���Wߏ���(	��ćξv��Λg[���ȱ%��>��RKR�y�H��%)�C��Û�R�ԫ=y�yQ�a�A�)�8�>q����޲�?u��dO���9���^���!��|�L^L�rl�D���&zg�.k䲶?m4r7�
6��L�s�<zP|��7l��OH�φg���U渍d�3�/O��](�� "/�Jҟ"N����������B��rH��w�Jr�1"m��ǕY��GLOI�F������;��F����n�c#�
X�yL
���WH/�#HGw~tN�������K�����(��\	K�~�\m�l�rƇ�2�Hw0�r�H�����2/3Wo*�y�G�n��Nu�3Zi�}R�xFcBDP���M��$܄��@� ���!�)��IRY5���Ivݴ�T��I�S�xF�Xt������KQJ|���&�(��(�(!�
}��M����a�����:�1����
��'�)k������?pn��i�!+N�S�=6��VU�G�y�F���eq���~�����%�  �����'?��Jn'��p��������|N�)R5Ba��J-�1���}��?��b�0����Y~1+s�*��r�����o���d���[]���<Y&_��j��+~gY'3?���aYL���5�S�?ȁ͋���8��{��������E)��ߴ:.����%��X����Iٲ`S�n=�6��J~���&q.&�oK�N\�V;�ʽZy��$jr4�ߙ�����%�d�חd�!
h�\��*c{�:�5��5�R�_sd�6�r����Q���]�v��U�tҘ3��3�BV8����׊��*l�+�Rԁ����*�V�U��,��@=�:��'��kɀHIs�)xa���J�q��L��ӌ$���4w��o\���%J��i0�=k������uDd.���		���#ÐQ\�h�iO3�i֑7���e_m�4�N�F8ܦ��^P���yA�� �db�Z��z���%<ptb�	�����t���֩��b�Ci��|�Fr�eZ�2�)�@k���D�eM1����w��V+���Y������O�$A��ܟ��FT�*�tQZ��!k;N��,��6�/>i}�t#�>@�d(��U?�F�PB��KYΊ��-��*�TI���毘�1���7�3ߕI���Έ#�N��C�*ݻ�mk/��4'5&�P�P�_ZY��.I=�5��F�(s&`�Ԥ�7.�~i�S�FNa��I�iO�V��ࠝ��d�E��X�&������~��U�rm38JO�q=H�}�̂Z�@� 1�8�'�R�+v�r�&�s�:�N��4��u�zݕ0��\-��Ւ�ŗ�v�g*���LZ���r(��J'[��C��}p�.G�����|w�4�ͩ#��K�qDӊN���m#>u�wPw�4����A�
Z�V�#�
ɤ�I=�Q:��m��v��Wc��=&���^ �����+1��C�Bmr�����T������,xo�5��(�zm+o���k0Z壻^m�'��$I�*>E�� q��S���1��EGu>�R�"'ɗ	��j��E�7����\o�2���yiI�7�w�y���G�}�7���א{�V������K��� 9�#��ka��n�Nҳ�:�|0��C�K(z��?5,(�`�S_�_�h��4��QgFmA��W�H��������7я��~�Z�H��?�8��Ʒ2�1x��I�m�4���V�@˘����e��<	(	 z\,r,�����>�H�b�׳l�ޯN�RyS�+L�a��`���H���"��$��$'�[���|*�w�΅��et;� eɜ;@Z_����c��*�h�+��u����i�P��NI�.@�F�4�E��c5�3�|�^G�.ԙ۱GG�\�]|�+	1���J��`��N�,�פ�����t�5�l{�h
Y���q^{N���5�&���҉�#K���#;z'2)23�n���2���9n�W�
��ߩ�À��8�d�
�B���p._�dK�k]*5���S[7�+2�?݁�M����I������ƹ&���˂)o�d.��Q�����ϩ����Ol��<�:  �דe���)O��i����ɾ�%�����	�a*��r��i1������R��M�q��j��z�~�X���%���Y�ߋ:
���;��]�5,ݵU��!��sY�QL���&TO�k�Kz\�$��Bn-���F���W���^'�Lu�c�;Q����O`�W'�^�s3wV�J�8@��ѐl�����,c����l�"�&le�o���-�	�1���LҠ`���/��	��J��^��R�h�o=+��%6�Mhx>�au?\�''��&[�8G4r���� @T��af�w1��`6��i�/�m�_%<�M",�L���V�tLvIU/]����䘸��1fܩ�-�5O�4���}�h�q�eA�� �F��J��V.�S�<5̋V�R�L���!Q�:�z��k�]��2tbk}y�հ
�c��W_C�s#�Q+$J�z+W�¦��J=���a�VP�qjLj��Ӣ�_l]L���4�L�<D�\��������F��#��x��ͭ��V�8]1��y�|�.�MS����K�N�:x'�8�z?q+��=�����C������iu�M�����G����X|I�<�È��k�m��z&Ћ������
l�M��v;���W
O���fP�	�n�"���䣴�a�"p�����O�z{���BH�L�t(j�Q��*�0�7>W�9�9� &F�nF:IA	D[,�*W��C��@G���ɂ9��)�_H�����qq���IU�?����4�Wٷ��J�,�4�G&��e��#FM�qA3Ho�'|�Xghv<��4�s�6��*%�!A@0�<@�-"�k��੾�<���$u�$��*v�K�"C���ht�XVS���%�w/�)g�(D�G9���2B�S��`f��d��ߡ��=�ź�����N�2A�IF�T�Sx��ۮ
�^ìV�QɓGU�A��ԓI���
��]'�d�����m%�p�ir����G���Ƽ���U�S��)�n�[]>�q�]�`2Z�j-C��?��g��?:5�:
�Z��w�!|yͻ|
�65ۮtC�{W`q�H�����y@�-���}U�X&(���J�3��m��Wy�2[�[�\>3��ń�i2�X���Wэ�`R���D�S�A���(�o�D��}��VwP NF��x1��\�GA
s��D�Tϳ��H8���O7������%̱�[��N���x�;���u�C1�� {U(����Vho��8�������8��w&˪�L�?0����h0ؙ:h�����}|��.ɇ�Y &���/O�HQLmE��/\��P�g���c����L�(�Q7�n|5�`����O���=~8�y_*�9H�l��c�N�*�=�װ�����@�KA��7��*
�W5����[_A�P,I�HQ�/��R��K4���pK������	�o����������6���p�&���G�Jx��d��j��iSZm�y�2�	����w{=�����@�颃�%9��廇�Gn�8�] �!l�����XS�
a�[>P�0coLB�~���N�a�ը�Q�R�	uR>��n2k�"ȘrΆ��ˌ8�o����a!�>^zX̗	�Q�w�
�eL<�מ�]t6��,.���נ�Ն�a�B?�ʠ�ͩ���hP�~_�����A�2��|���<wbN1� �gVa��;!	��p\TKJ���S������� [���d�}=�~�l7��0ch���צ��&���s=w��;
�.���e�n�u�Pn�!����m�h�(��6�z)�5����������T�m|�Vh'�{B̣&� #Rq6|�6�2�S���hs�U+�%}�����1���@���d��b�ԈT��J�p�Q�w��w�^4��-܂�ZVg�G�ݟ?��
O��t��䇾S�t�͔���d������@�DAٖ��`"c[�`T�Õ�;�����wq��9�*�PV�Ɵ��P��!_3_�l1�%�'Cc���_n�Ł$�n��ƛ���f�R��,:o;�S�R#v�Γ5&��$�T+�)ì�����,Yn����j��1���2�b��<��;�����4:N��+�m�
O���ݖ��<ir3�7B�;�t�3����2�����SQ$��7nvS���̡��J�oV����>D�B�[=l��~�,'�~����.���T����E���pC�o����_��sB �V�|D<�{����`�����|�����Xa&8�ɋO����4Ƕw��F;..($��.���l	�t𪎮�bP:!�\�"񖀯3����#��c�[�ye%��ߘ��bWM�&5���I�6;�H癛���U�@���H�prz������)�A�T���� ��FxIsȼe��l���Qϸ������t0��FR@Y^E(b���h��o��1���m��qC9}�_o�����������B�W؇�Q���nH��/@B�o��8�������l����z��K�s�S�<I����[X�Zv?��>$��b�>j8}G	Pϵ����8�����C3c,�� ts0a�PrZ\��5N��8���ᑩ�]y�v/0��&O����p�co���T�*�5�����d�躰�GK�0HNF�[(C��X)i�e���(x��˺�ȟ^���Կ���0ԥd�ǒ�7��j����/�o�F��
N��s�y�}@w����W���� + �TL�|K��=�59��ɡ��,���&�:�����D�%?�9�K`�`�)iu�2���^2>�5����D������%jW��{*��²��{���)�5�b��)��|=0O��U�ı�}e��"T�Q���Na?�`S��}p.�ilbZL-ɿu�Kܽ����,#�\�!��������=L%���~JǢ�y��� ;xw 9xfz'cv4T�%���	��%-%����RE8�Qy-�� ���>2�L:G��E\N���5PP���Τ,���D��s��.1R3_���iXG��-���,P˅3{O����F�Ö�X���<t��F�lO@A�U҃�Y;�U�x��tMl��-���J>mQ�����Gү�f�# ��`v����%�,,J'�=�)�A��yZg�}��;\,*��*05)b���|`��Bs����PҐ�.Nɣ�I��j�/�"�Uc�㗾�h��`�	��_Ǚ���x�#�-������n�W��j�j�d�@�|j��nWp��Wsf�mFM��De�&J�K�-د�(�|��N��_�ѿ�>�� ���]��̭E�D
��ˌ��� &��#r��ŃY�U�Q��۶d5Y`����u� ��������"��V2�8k��&[{=-Ŝ��Է�'�0Iy�l+�����4��w'{���k&��u���F';h��_y+:*����D����
��;Qv��)��1���vV�R���|W���$Ѥ_B�f(��6���[] �{s���:�`$Y!]��zO�9\��dѣbF��f�Z>�ה#��l4��.�J!�I��m�� ]=/a��&.*z�B*�򩿶�;��JI�j�s�I��k,R�e�3�|(�^�vրqŹ15���z�v͜��sc	9�tN�|���5�8l5RsP{	]l���{
c���b<()�1�����w3��$:|���ғzσ̑��dE�mFӾ��Y^X��ٟ����\�`�vT�~#���s��}����}�ьYAZ�`h�r�����I�K��o	p�?AnO	�cBe
x�f-}A��F����m��l���qɣB���݉�z26��	�������1A�vL���R_ˉN(/IG4t��zT��#�`~J���f_�z��	]f��Y~����C��Z(�qHAJg�\a���GdU���)+�Ly)��Xl�p�νDo58��I~��7��PR���>��Hy�����P���ׯ_؆V�@���=�'՛ ��y�j�YoHz��� D"J����w�6��=l���UL�(�]��#?T4]̺$�xN�<�k8D ��ĸF�#��>��-�!�&�9�~�f�ݾ�2��1�{��2��⼒ ]�5�����8��*�S?�SjM�cxj�T���Q��Oz��c��E��u�+�AY�ͮ�|y��O=��*=�0ێ���"h_�RN]�&�#��^U�P�,5b�qj ���2�R+0��VY�)����7��%�������bj ��p^��g-Dq
@[S���aɑ��u'Q�U��f{�8��qK6"�u�}�d!R�Q� �P%��L����I���9�ԉ|�h�6���7]7a�~}=����g���'�^8k�t�m�+ֺ�!:�>�K����[�5����-,�2t�r�ppԶ�%x�M�[�2�E�W-�P����sz'{��n6����	��x{^��C������X<m�#�z&���٨T�_Zρy�3��s��"�Um,��z)�����J����pC����py��F�X��V$;�{6�5��3?��Q0K�]����c=^�ܶ�W��t�D�d�W�
�^nw�+s5Ft��K+a4s����%��̦/Su��Ns�cLx"Y]/1L��ٚ��d��< TXV���:�3�{lqgu�	��n`�)�K�V�g��|�&kqQ���u*�0�wO��t� ��`RA��0,�2�kow�~�w�l\B���_#?��8��k��F�5m�8��.p��pK�zjm��c�����#Y1����X�����C�����"0����D�f�p����I��c,U�{�gx'ܒ!��?J�0Qb'I�����8c��e��1{�~�$mQ9t�')�a�?c|�mm�~b��gdR.�/	��4�d�v� 1u����G���De��ܙ������#w�X�㻹-l�T��x��D�վ�/�Z�nN��h^4����|+��ʲ;؍��E6'"9nq�d���g���EQh�}
���t����MO�ݨ��O�j`$��b���}��V�^i��k Jj�����A�\8@)�[�m�p<f�2���!r�.�M�\@� ��P:��u t �}�w��3��z3^�?���u=K=���rĶα��p1v��k�V�B���B�g�� 5��&C'	r/P���VL�TGpJT�8�o��aP܀4�
��+�n��ݨ9��z�F�\8����rOL#���)=?}�&2v��V�M�[g���m���1I������4ב�-�(+R�>�,����G����Ԣ:vB/���1�O2�<]�j�F.�����H��Uk�2`����6���>���D�c�P	-��3���a�Z�4�J[ļ����
2�9��� �O�G2v�"�X�B�a ��Pꈌ(4�Vo���n���hO.\/&r7� Ib  �v����μ�r�`�Z����O��
���������=����������RvzkM3�l�Ƈ��^�����5�ʄ��D�Z�U �J�o<��*
�9��H��Lr����J��\өx��P�*����3p��j�ّ<���
'�KDݡ�"p������K���5��WQ&$km��v�h�fI�/�$Z�K!C������ 7�t��f�9ؑĚ����,
�1f�R�)�B�v�A��tl]��c����$|��?�k���{#�z��$X���	#f^"ƾՎ��9����W�v�5��m��L/�`��]�F�-`��A�5�/T�-��ņ��|�8[�����2r��aG� Y�hʄ��!��q�:#����+�l�m9�M	JH�b�i����[����$��s�Ҧ `���)X����2����O��ܴm*A֢�~�ld���x��cn�G���g9��ǜja�7�O2G��c)p���%�F��5u�o<��#v͊N�����D	&�H����L+}AҪO�q���]�܅�	*r`<$�T5ֈ�L�5�C7�?�VG���Ǿ;"������nUM~˯Z���r�8+����C��N�p �H��-w�"��Ivl!+s,��6�(� ���s���w	�Ū[-�K��)�I����{ٰX��-���\�~d0 	�U��<������r0�M��r�6��X;Vq����0_��?`��?~�vʆ�
rL�
J�%7��׳�z��l�lԩO���M=�_�;��<�f'!����J6��[zd��*{���7��,b^[3]��DJ����ŷ��w���,�nğ�.�+��f��m��<һF`��z�􅲉�Y�:�|�����56<��K�S�%s�EqC^$��7��lO�|M2�_D�w������{��3N�h;:Ɛg��x^�5 ���X�@X.�k��j�D}ڱ�&�pv�����`=��|H/G{�S���`O���V�h�������k�?���ܗ�����Q���]e�kfR��М�|R6J���w�a��>k��D�*�����g��]�rP(�;�A^�`&搛�3K�L��;\�ov1���[�u���>e�-�R=L��M��v��OQ�x�ji��B%�ht�4����S�{$9b�R�E�)$:,�ëe�zt�ÏhK���Q�&�Q�խh��OUUk�C�C�r��s?��|���-�����*���ʬ��U?i 7��|f=)�2�g���`��R>{�+��Oʕ譨Ogn顶OBp1"���5�e���1�vA��'�v�F�%�\k)��WN������<������-��]��D���0��n.J���>c��Ѱ�\z��%���+�I�w�����Vgv��ژ��n<ܰl�$��vZ���&!X�OK_s�^�*m�`lQ!�����F��Ȟ�
�9Ȑ��?�$�yw���x~�F��$j�=��&�p����5iV`rt͓!:�������Y�nyPݎP
����ӿ��-�:��W�a��	����Iț� �(�A?�q��=��tP�=��pĩ��K�dW�ǯYW���K'�V�Nj�r/#R@/��^OG�=�J(C�w�.�/]�y� �){_��pL�f��X�;��R���,�0��,���H��.ͺvt��Ht�!��-�A�(�d'24#�� �}I����v�E.&����9PKu��$s��>}HQ��Ҝ���M�ʙa�N!&���,��4��Q��D*o��^#��A�@�s��Qޣ��ӫ�w� y_����mh����?��9�Kg�eZ��J ބ�����qfIs�%%>9��dyL���A��R����jv�c��lŃ�C�.x�"�̥�������x������r������!�0�q�]���a�S����7\kW�U�]��¹C�s����9!g�	y�
~�,,��W�x�� �MY��N�z��{����>�D���p���k��OYo��O���<����W�P$�fka�q�Y�������F
Ե5w;�|�	�"<������Rؔ�o�n�.v'o���
��P�j4x�[m�.����[I�{�e����A�g}k��de�%��5�	��SH��5�� �Hw.?K��?cfXN�q��DGHjf���8��E�1N�rߊ/t�O�RH�rK�fD�m��DʛͩPX���LiQ��&��f�_���R��=�6~�"�qp&ֿ�I�X�3Uȗi��;*��0��� �3�$F�RS%�P��N�������>y��8И�D5/OG�:6I,��uֲCItq�^7a�$[?��~��r�Fr`�,qWߠ����&�z�-{�"H\�=fl��(F����.�߃h>j���?����V�͒ZV-�C=Α��?�қ+J�,wI�>���f1��P������!�W)�_��tGᑂ>l~�M��k�x��Q��t��s�MC.W6�k����Z�qGe����Ɗ���uӰ���2W0q�|���:袞��+�M֧$Y�_D��B��Ә����P-�+�7�{��Mk��YTI�����D�X�͒�h�	�|�Q�f$U�?�9���� C�PnO@Kk�+��/fc��ʠ1���md�����0��%���&b͊��GD :�L�IZ�~�;(MZ�r�Ik��N�ѡ� ����|���Ym���� ��Q�е�/�
Z��u�fC84�Ac��kd�V޵j��c�<ц�O��-?NRCd巋�-{���oeU�`���al�>�0W�[�H,[D�xJ���[��Y݂�e�m�Zp*[a�BEM.G3#�$}��Vf@N��L1���}݉���F�E��gø4�����n�LU.E?f�Y�u��� T��x���;�������J\RO�lA��̾U�,1	9N�6�� ���RIٜtwq�$��%�%�Y7���z�
�=��HHD:�C�ֶ)	��kwt������e,�ȡ���t4�V��34�`���pL���B}�g� �aބ������A����I]ߦ�����+zl06#�pr��c��䞄zߡ�{�ӳ��t'R"��Ԛ_�Z�8_ŢAGrc�eqOJ�nI���_��Uxc�p���M�i�v#�)��Y �S�&)(�= 3����pLh1(l��$e�V������{+�(O6�"-~�B��"���⫪�q�ס(�ט@�4a��Ԧ�}���Z1� N��0�]p0	�L�G����L����kD��
�$������ŹKl�D���prڮv�y��xW������fZX�J��^x�`d��˙���S�"Zޫ�>g�㐯��5$�fH!�����^�~�.�-���Z�i��O3u�9��y�d��#Oͽ	�*I���$�˪�W�>�J/[BWD`=ӻ��x<Snu�����H���V�^:��g���%h����#@V�YO�	�~�9ʊ���X�Hi��R�IGo��N� �Y�v�؝��a���G�`��h��I>��%�OR��[}�������A`jw��VvT>�s����$z	��@	���:ޗiP~W�V-4�Q�٘/�3��q��J<�<�D��� a���*!�
I�~I,m�<m�n,pM���'м�Ƀ���o��������kyK�U�ͷNt�Gt���d��oJ"�w2}nل�O�E���(�%�3��%����&��u����)"�b����hl0eR�0F��@=�?��}�^^g+; �=V��q|yx7�'W�i��ʈy��A�w����D6�Cql�m�'��|W�t��u��,D1ma��5bø\���]8Js��&;�P�ƽ���(�[.��@��x1k�&�lD��c��:^�bY&o�]����db���:�݇yD��*h�_�N}~�hW�i�*�W\����	Őg���I�Ǘ&?�H�V?l�=�Bk��Iq�\�MU0n�_����<S	��m���dfB��F��m� ��\���D�*ca�V�X�c�O��˫���|�t��;�s@
x�K\�Ma|"WQ�L�N�)9[�t�);uܓ����)yD@w	��[���y�&�\��W�/��9��R������3Z:��T��M[���_�t\��,�.�!Eɨ�^g���Bi���1���/g�)���(�!��V3�_����dB�|�ϋ3h%�DD������r}e-�"	@2����\ڃ�7.�8/e>�"∁�2�(� )s��jH���O0B�4�q��ӫ���u�儌J��Jr��w6��{n�&��v2��Z��cy��L����kU�	�ޖa���5	ܾ�ހuPf4��%Zc�{3�yQ �rgi�\���3bS����r�����IXI���c��܇�d9L>\�=�&B"�U�4Q��&��rP�@�	C0̜g���n�&��_|��a*_�ʬl(O/x$�i�ko�"b���J���`��n��ކr$s)�����5ܹ�5�iH2�f.$�L�$�H0�����?N��y�J\r�#�H1ċ�����M������k�3�%���LK�G;gk�j2�$!,I|�F�s�g����`��+�^fG����<��b �_���f��U`���z��`V��(�����#�p.�\�nN����a/�d&��]g��h&�b�^��ZR�Nܝ�H��}���*|PVe�t��=�kZ���P�Ăn�X��q�!��heSF�j�s��hY��hI*�h�m��ų� �Z�eB��e�!"�D�qb���U?�/�4�	�����
U`d���S,����O�H4��� ��*F�zU�vַ#gR��DY	^D�!Rˤc	㺸��֌�ߑ��3$�Yu��� �~�N��7�0jm��G��6�E����5�~�&��M��R&��]�����G��S�^y�[(Mk8Kr��KԢ�xL�J�����x< �N�n��^]��&��.�J*lrd3�VeO�R,}%����a%��F��o����藇�
��Jg?����ܳ;0�>�0�;�5��a�I�Z�^�-�T%����M:<�3{��C
�6��2�����T�YG��H�1��\uR��K2�)���n��?���0BYLc¨������VΊ����.v_��)�ڂu�W��  ;�ȼҾ�<�PWMf�n�l��K'����~���'L��UF�QC11XI�wѢ2H�4o 2�?"�]~J_�h����P�-����5� �����&^�ȶ�J`��
ԔJ�9�+�m�`�so���D 3���2b��87�@���x�����3������*��PCYN�~-��e�!�5<�T�5����,�Q��H`U�X)�FIJw��K'�y����rj@�� zm_(��U��q
�,Ժ�i=���u�	~1T��E��Z�*Z,�?��℈�t��p�j<����0f,������\<7�c������:��[]Z�-u�yIj���� ��I�&��,/t��6Qa����ڂ�M�[Ou������B�+��g���h9=i�S�ZC/���c��!iߕ�^�>�Z��c�?��g�͆�"8��~�����J�9�8�:�1��eD'��B��^�M�T\{�΀u���`s
k��(�dE��@�*�c�3b�8^�5ŔA
�η"��#��t9o���K~	x�v��3��	'!��M����Ꮡ���K�/h�QAm��S/�V����g��U�6�2еQ߹�,]�U�곋;з4��
uM��rLR��D��^��;"YU��\sFֳ������I]����F%�*�:��$���R�N%-���  Z�����Q��Z��r�z���Ă��<&x�сe��1>'�hu�����J³ D=?ħ&3T1wz��m��
	l*��`��aA@���DU�(���4qg�/�:�J��KD/,�𩧳�Q�\��6�5F&����y���"y�
�*m=��պ1KG�C��܏�C;�:c�c��#(��϶y�YR+��J4�;���C0IAd�!����nxҍ+J23⪑�N�;��ϰq:�S�8dC/|	��i-!��,�jr�e1�4�*�U&q���ǟ;k�� 2�fUr2���,\���\�p���U7���;~[AHӸ �q2��-69�i��1?�ƈ";���7�#���D�G3{puS�
�@�}G�A�^˹#����j$��McF/Wv�.Tc
�_C�t�m*�4�t,2��>��ϥ���	�+��{`�P"�C��ׇq8���-�~�[����;"h�cal���C)m:S��uk���iWL<�=6�=(˕L�kM)6���eR��Q����.BȆҫ/�M���Fܾ?�p�$>��M��qf��5�6�>���)���/&-{6���ĜcŒu�!�uI�p���U��Wn�Az�����n���M�x���Rc��/K��8yU_1w}���)��4�ui�v�F>��
$1����y���?"��i�@Vae�fF&>�ʮ��LU�o���)��s�=�%�Z|�/�G����갤��y�L�>R<���51(�YD	��}2���sM�پK�ӧ�ҹi�A֜ �I�ݦ��|�q#���]�(4�]�;t;��A:���Jn�i��ޔ�©�^��x.]�{2]fa=���6.`E-��^@`���\�v+M~_�;���o�#(Z�~��f�#I���V�l=�u]\�U�u1�?k����`���$%S���} �y�&;$��8j��(���`�Ww����&?����C~�Y��J~Q2�9;嘵��b�����0X���b"E��Ê��!�QR�g��_����eT���ξ[���zAc��7�1����Mԯ%eR�f�'<�#3ʟ @I���k@���H�&����'Dن��dj���:Tj�֨���e$L�F�� �����*�LLr��9���1����zc@�w-���KD� �# �PI>�^*�z � ��CÓ^Į�k`��5�� ߐ�/�sݼ���%�E���jB��擬�#A�D��Z�j��b�k᧺<	 �/&cFu������!.v�\�>�����v���8�$/uf�Rlv+a�mʻ6\���a�@,Ҍ��0�u
�:w����{���D�_�}i��@�t7�f����j���l^7���Ԃ�I���ŐE��a�ˍ��P�x2�w�aԥ�
\@X��&����<��+�本����?����+������K�)���33v�Bδbv�VB㬢Jd��to�C(��!U2b���q��LA�<x�s��
~o�� d#$���:�6H�������ә�z�3�$x3/~�w�#b4��c���<p����\�,�PT�+�롙�0X�nr��)�k�W6�:�5�W�jxs�j�gVNn|�x�.���71��9$T��$��S#}E�m?�i]��$����۟w>E|�ת�!���ꎤ�O���І���Ψ+���G�BVw�]T�m�1�?�m['4���6^�{0�l�n�|���p��)?��Y�>��E��h�Ft�]t��g)I�h�0���TVT0@�f	Z�v�X]V~�P����[�݀�&����7����o�<���:�H���T�x�+P�h�˹e�Xro��c�a��^�5B�>\	!��}0l����H�)��  �U���lIïǧ9OQ�I}4��PQG��h��z��s���P�M��6�o�+��q*���g��+ׇS{]��шeE��bp�涔���.q��{d��Y	��`��iVŤ�s1\q���E��5�1���_lJ��ӥh\����_���)f�M��$8e���N���=+���_�w��H��+���9ȶ�]��U!ߔ#2��7��l���TQ�T'����Gg)q����Z%R�8]��4��ehkv+���6G�
�	��&@�7��LB�I�_����?ٟ�+����+��Bv���R\��P*�
U�#TTcܤ�%$-h�Z;�	W��a���7�w�
'sn�jbt���8~έ�l����.�Qxd85�K�A/��Cy�;���֪@W�h��%��/bܖ���Hi�}�;�,���P"L�}(o�i��|(�x����z 1�g�K��z[8.��ua��˜i�k)sqn���l�z�'C9� ��Ns��A�0O%*f9���Pm��H[O�@�\��yI�ħf�;�!wX��_�N�����.��p�3��o�V�&�B�s�E�\�_��>��F~cևe�.5����C�pQ�.8$v`�Y��4t�����I�#�������,��A�I��pg'�g�+]��5����kh&��8ڱT�����BV��:W|t/p\{R�D!���a\8�� ���v%N n������y����G��h��%�"Y�ʹ�TB6� 8C&�U8�˜��t �I�\�qS���3op�'T��-놴��$8��us��l]?T��x�Boa�����T��ȟZԎ8�vf�����'����t��8Ymcq�!�H�
6�*{gkĭ07yE������o�.�
q�ֈ��Z,T�����E���������^�1�{栦T�!���5����o:��X3C9�>���0�=��\��]�B,@G���aJ,ӈ�")�]���\�V�D��s��&��	G� =n$6�4����4�KɁc7|n��S��U^���^��i�N��._f�|2� ?��	�^ݯm���l�Gg9��9M
L��0K�<>�D\İ,hHcV$�ɉ_�23��R;	���:0���݅��Ӏ��w��ӛ���9��db��� (UQpc�z�^
�J����n��e��ZpZR�/Vׁ��vG�Ն�@�� ��%5��u^�}�ϟ���>�*�M��O����%����_*�-)��[�	v/�9*����k�s�'A�D擬+��G�r	��q`��7V��Nu9,y�(�W�\�U#��w�^>G$���$tk�ĝ�
��#��d�]�k�������O�cO�ǒɎ�ݙ��3O*C7��K��Di��ƀ.��D O�d�ϡ&��Խ�x��g={B�W��52�%�'n���{P��+��e)"}�X_7IQ�R1���7q]$ݓ�h� ^#&�%��s��3Jc%x6Wu�����i���K:��h���X�X����׶Ѥ���@�N�he��Q�_� ��2��@�F:�I�(��p�<�.�� ]����ToE�g�F������t�g���.{{4U��\��q��4gM�t,���1�x������R�$$� p�h9����#��].�'K��Ft�G�!����,��mT�;0 �wS��AI�TB���L�~�ba5^�l�@tg{�to&f��ʔ̞�i�C�'Y:'�i��W���`O$L&���ř�_�r:5���k4@P���҉5�bW	�K��$�7E�u_ŵ�`�TvR�<.�o}�.��U�vsA�{k�$%fT�fCP��u��?
����r�N��Cz�"��r�Q���mw�dY��}���/��9 �P�:����{���j��\NhN���h,qZ0�]~��K��I*�i?W!���bĎm�B_�D;Q2��<�"����
�!��gʾ6V��_��!�����g�?�tJ}� �q�!L�/��܎��v1�������mǾ�� Q�BO�A�M��]13]�uG��p��=�K�8�� �#Q�B�٭����f]��	#�KA逍��� F�V!y	��+��ɥ����~���i�mC)D9~0��m��W�8�}0���n��/KYU.q4���޺S]�>�����{��Q�`Y�ã�VwV�q��R`��i�/>��p��Q�m��a'�_���r���]��g.S>�b]1��$"\]�{G�i9�}��6n�;*�~�|�����;r=���)� jw��z��L���{��Ú��w���w�h���,9�}:aZ<�S��~�Vͅ��\^�ZT��Mȱ�w�j�#��I��]��Yв(��s��s��+�%Z����P"t��<���Y�X?;��@���E���)H0*�+�^�e5�j�
z��6�c��2�#Aí�iA����S���z)�ސ$�N�Q�S��X�'�v' �����/w�n	�C3�z��wF`��_�}X��-�_6.��WNG�f:��ß�����=ݿ�DH��d�<����*�=EK�@̟b�C��+I����Ivh���m����Ŋ���B0c��C�v_��-���8��kd�7���i�9[���!��cx��@�˰�%����t���qˮ�S��̷
�%cMVQF��&l�u�8�~��v�>>g�B��K@9���_�������t?`��iqmv�qZ�Aɾ�����!�C(�N��e��r��ӫi��g��