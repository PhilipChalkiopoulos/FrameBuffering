��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW��'�mҳ�۫xv�<��
�5O���q��z*�\�"�ł}ʙF[BT�8����f���Qq��A�?kQ����#���pN^�}�2P��3�;��UD��UVҪ����7�5G��Ξ@� �Nn��=��w�:���"%~*�#��Ok�����N�S5=������3֬j������K�/����9����d��B��}L�d���[
ם���Z��}����Ϧ���h�8�������&(�uv��-���T��8�,��O��ܤ�o;_�m�d�[hȩn�u\������J�([{ s/�H7�"g�>�4JhY�KA�7�~
s��뗗5Ѩ�KO;�АA���m�����T���?)bs���HMvp��b�3U�V�*�v���/�x��qi�ZR@���-�e����{�&�`�5�B�"���5���[xp�+b~w5�;.9�)����!�u�u�7^�N�ۧA�Wa�>,��h�g�p��dȨq�Q9=[S:�y%���Ó3Z�	�ZZ����$���:��.2�`ϐܕ\�>m6��|i�І|v��5G��TnB7�k�E_��\�N��!Yj
/0�I����}���1������U)��fQ������ 	���%��5�DI��Э���ݕ��u�Ū��ɉ�j��'"��h�M��$�D����,+���-�x�Vߠ���cH������a�v�Ӛ��0��UT�/k��И�:8��5D/8\[S*�rT@[�8�~�V�V���Tp���� ��&W��^�eX�G��<4XIO�����Y[�O�b��yJP;׵Ӳ�$�"��λ�8���3>�\�U�)Yr=�O|��O�<n+y�j�Uo:�E� :!��Ҙո��F�A�P�ژ������Ȩ��g���d��#فmU�Q��z�f}�ϥ��kJ� L4�,R�:%����(F�0�|�@�\"�-��xƦ�w�xz�	p=��ŕ��׶�zm_@��賜�?�;g�ܫ哩5p���JG.
�&��%�L����[��'<~��&�aK��J�7p�D���m\�T��*�藩�?��Z���R�8c�,y�DS8S�f��?�,9K���4x��4Mg9�o3x��IXp'���\�����sK�x�hZ�D�����x�r��g�G� fp�}B�(N*��"d�����!�=tB(q���3��=3\҃>X%�J��b�Zif(Y�����o��X�ջF3�AZ9G}�(�7�[��ҠU���\�Sc����G����K��>)-i���3��j���S������N�'�r��� �_�]�a?�X` V �K�(�B�z�ä�Gm|�{؏�?6@wPUة����Q8��D'l�Ch��՛l�������B�k{��3�{���q��3t�#������ �P��˗�6EB�"�}��Z�(�H�֋ڨٷ��M#��[�l�����vo���s�`����oc�L5�\����ť�>����ݯ���j��-��`Vָ�_�hlA���r�Q�K8���T[��R�k�Us9��!!��B�&UK5�+���0NP�W�fb�gXx����{C�t&�F%�� ��l��N6.h�F!��0�qC�����Ь#!�|���E\�/�I7�<`I��{n��o$}?�7m�E2ƙHOm�����(���A]pTk�]�ue#~��ty�t�N�Z�a��jt�ͭ���/�E����6��,���
�p�A컽��0%�,j���I;ga�Z����B�ו�}��D�+�h)��e�n��M�Z`� x�a*�YТ�)"��r���33���\���|�Z�r�E5 Ώ~ ̖�^�}���)�33䙸m�Kq.�b�4���-ՁX�X�UL�����KHG�,��}U��k!=�	�}2eD2��c(�D5J*�<t���|^�`7��L�bъ[��"��%���(�o"d��Mfe>�iL�@�8 l*���jG��󯇿�������o���b��;j�8�u�A�_d2hc�k���<s�S�l#�A��?�P��T����A���`�\�*F�6+�z!x�r`�=O1 ������������|R�3f���K����Fw��t����i�
�ŏ�A������� �@�to��e��ܶ���lm �����iU8�*��?f7�܀f}����^Te��G��	��{��,�E���b��s�e�e�S,����/�/NY/��(���	�GPE��l1�Q��1.F$�'w�,��Ņ}[��*��Y0=h��s���Z(I�4C��^ �(y��eA=v
Ѯ��<1�=-��:T�T7�+�#�z����iK0��3W�З99J�����Y7Q��s럢HI���a8�[�n�'��h�V�^���г n�}�K��}�͠B�� %;Zm�`ۥz�!�o NH&��6�:~�p:�" ��i���H�峷�u�a�rw6VhP�Y�p��*Qq��@hxStT�a�J�����0�0���Jf�����F���OĲ���t߬�$q�̄�AO9_fn�/�hQx�[�v�ɍԼ�n@�<�H�)P��Z��	�T��C��G���xµ���ˎ��}��fz]:�1Qު�Mc�n���=q���5b�P����)x+�<�@eu��o��D�5�ddᎋ|��t�[�[+=-��d����{�?���I��c%�X.�-�|b�|`Q��ά�1�w��D�KS5�#Dd�����W���6�q��jf��8�^��m�E������B�ut�(��o�������<����r��xAy���Ȋ�=zD̴�E�N[^�i�ɨ�Cdŗ�`�������K��iT<h?ǁ�+́��] �l�L�ҫ�;�tn}Ry>��!����#T#�"�|��Ti����C���,��j�ʯ���-�Rp��|bI�M�k�a���	�h��T m���^��'��Dw˲p�1ѣ-�s}{�P�k���K�奁�?���g҇71��S�2m���߭��=�O��6�@�R��:�P�s�D��Rƚ���9ʜ%�w!����J����.>z��|p�*�+�S�K�9iV'R�0;�2SL��v;�����P7M�(��R�Q��iO��nI��J�D.�q��q�`5����xO��o�kS����l�MFjx\b����H헢i4��ʞ
F(i��=��r���;I�eg�h�:�lI|����<:���2�'��ׯ안>�UO����C尲��#/��\�oO�����`\���U�Ȅ����LM���/���d��FP ��T�	W�k�b���d�uml2�����S��)������;�a�kFlYu�M�ajrZ�'�G�l�7����W4uΣ��F.x��������W2S�;�v!��';�݂�/|�O49B�����u�/[�gO�>Ap=0u����$+}��z��ZN{,��=�q�4�<z�܄}�2��Ī�B��#�hu^Cs��Uq^]��ӛJ�t�Sr���N$��%"�wx���}�Sдq.� /-Bm�K`v�3L����
�BI.&��Q�̓H��Aeئ>���Hp��w�w�}z�9�f�>@}d&v@9IM�p����3�	�"�ƌ�c
�]^G����vB�wI!�:ƴs�2�����s�1e�&g���HN�t�@�/�?m�x%�s ���V;�_�﹪���B}��̝�KٙOٌ� OA��g:�Vu��*�/������T2�J�"�����Q3!8��Eqae����kK��j�sSZ�&݃�����S���|N�4hX����#dCb]��a�@6�	m�V,�
�n  cA�%��0����4�wWKI�Iz���kdJ�����y1�Ϲ�H�?i��z��#�S:�~z1|��tk��ޔ;�++�X$.N��'�u�V������`��`k��d���f���C�x2v7�^��j��7'$�A�Ij`�*W	���M�3�;������tV�*�:$,��v&U}@��F	j����Gv����u���+�gk��I�"�h�ӂ�+��C[7��ԡi�!Mpt7�S��܆�U�䄞Ç;tt�!��(��Km���{��K�:�������Aļ�}�Z� ھ%^�x[�^���b�q/�"mc'�d<;�J�q&��ح��r�`��c�������֐�'p�ZV���U�2�h�ɽ���d*��}�~1���
2�P�<�z��&���4���:�c���Ϙ����������Iׯ��9ϳד�s�ie��������f?���p���|\|JQJ�ۅ��	"��קM:��2���L-.c�{3yP:؛ԯP���Y��[$͹�r	�O��� �%v�N>˟!R�P��r�yh�7��-�µN�>�����#�R���"nƩ��Poz�h���CQ��:p��L3��!��
�8,������T�Z��$��-�H�~�ȷ�7�8��P�;.�$���|�ۺ!�A����������P��Ų�\-���0�z���{j2��]$�L�TԲ>��b�����]NX����ŭ���^o�K!+K�R@D	��B=����ÿ�|0|aUAeisjc�1�\� �7�����8#^u[�j\�w��c%��-�4��� f�Ar�k��U�wF*����n��M#�N���١���]^+�nHJw�X��x(�����d�G6W)N}���V^׿�If���mT8[�-���&��� �j!B�W��+!_�45�E99s��Q��� �
�T��A:�^��[@��Ɏl9;%�p8`��ڡ�?4d��@�ՏT���%�D?���-�����¬u���RYa�x�I.�S�Aw�;�e�zфmK�6��4H�2t�ET%���:��hr��ɮkB�{*�;|��E߲ɨH�B7�����i����K�ǁ��7ES�ૉh�TE f�AO��=����b6O-ٟ��z"D���ߘc��˼�������$<��pڕ%�`��Wde�4�
�t)��
�m�0��8rTE�#�����:�7\��WF,�)��E"��2i�^Fι�<F��5�[�����m��Ps���4���}N���J;��𥸅I�»U��q��h�"42�%��F&�p��Z��Dc^I*9�m���gE=㚚`�J��*��gL�6��t��M��UR H��K��5��l�}�����
[���6Q#��U2�D�	�̢�o�n�@*oսr��)�zΎ%�7a�j�Tl�4���m܋�]M+�"n.��!��Wb�0y��`�@;=��g��Be����s�/X50�۰��b�O�f��������X��:\ �wIN
�A��u���Gh�B&�� a�/�Bt[����ɘ߃D�O���KU��NC��
����ȯ	�nowc��C�g���2���*��]�tydmx�k^�n���\�]�8��O�i����.b�c�ހ\̵����C���~���Ƃ|�B1�����g(kH��S�R$��w۬|��oPST���`�78-q��,��j=�yL-�03��52�V �nO�D+zO!�6�?�S?�$�n�v����h�Xx֚S�V?�Okz1�^��X��4\�h`�(���,h^IP�_s+7�V�`��IZ6�M+��!��6i �����9�Pҭ��*�G��A����5i�5?臞٣�;��3`u�qȫ:|V��_��.@X��V�a���ʩ���]�F�EwI$!W�~�dn ���Y����>�k٠��Y|�4��8��F���
Z�(��J���F�u��~ִ��
c�]e��t�챀��,k���GR�w�e�y�=m��ұ��}ɵ%m]��`i3���~�_-
�Fb���%{"�%�)�zrc:)5}�@+0�O�<s��YEf_d�@��i�ø�Y/�vr[Z��I�Q�����-#�̑.�r<wm1��e�X���ViA8�I�}@����M�� B��CZ���R��%4e����M���c/|��υD�r�q�i^̓X ���fc2-�O��Dd���Q�/Zʚ.C�@yF�m!}R�;���:�ݢ���\ї�ؿIߚ��}ȗ!�3Q$V��j��,�Xp�I�y@�M	&�dZ�J�)���t�����o���xB��/qP/�oLu"�=M�U}Cn��u��6w��n7�3�g�����+r�kd�8 ��Ȗv����9�C�CdQo�$I9�#�xw�=:<���v%�� ��ʵ�~ȤdO<�0z��+�F��@v�p!���
y�?9Y���c, �P�Pd�F1-'[�T�����9��5��i=���F���YV��i
ɵ�#�)E4��C�������>9�tO�{tsZ��SA"���
��2H��X]���>gZAq!��:Cd��i���N3��7����{�_'0j$��J:;�k�H|B�\H�xr��&zd��бY5:\6��b�z��V[�* �M�O*�L� U��F;k�2=�Y��n�_�U;
\�^�I����?��{�ק��n��gJ@�KZo�{���!սE}��fE��fp�,UQ�.w��_����}�	C�oW�*�*x,�2?N����Qd��v�Ϩ�Z��?ʘޥ3
��a NT��ǭ�ǩB�`�Ziw��ze	�"8T���k)�˷c��9WW����;��?:_��o��������W�O�6Z$��B� �Ɗp��V�x�-) ���#ɣ]:�И��L����\4�`Uz������s!jg�u��r������\q�H'AԷi/���JdyJ��Xy��h��u���L\�����?�;[=��jR�3��h˃�P��F�~=��k=8d�Ay�Ua�bd��pC�CW�e�#<G�0]�n�A�0B�ɒ8�$ͤR��΃�{7���-��辣�>h���	=�����E�$Sم�����V�!���D���G��k������Z؁pT�6�=IO��ч��R�i�`��!b��]W�v�8E�,L;鯌�k;r���j�H7y�O�&�[����	����[VNýB*bdl�e#]&�>r��#w�v&�����b���JtM��둄Σ��tV��;�_ُ��"E�]�/ƚV��?��h�T�?}-j��!y˙�M� �u�6��c�~�:>��b�d[�۬=��Qǜ'we��|�N҄f�}�Z�W'~�s��c��#�⫔H��y�|s�����*�휎7��i/"K�P[H0�c���쬰Of1\�̶'5&3{.]�Lb���u�
VFKI���[��O�t��
���� �*IC
}b�}!���3���.u�|A;?�թ-���������6-L6^�W�{�.�ʕ*j�e�)d",�"�J�!����,��K�	r9!�⽰�B��_W�G�K3d��7���a���Ő>���ʸ���TI�K�q�(oC�W� ��)�RݕfqUiJ5,hKئ��H�"XT$�K�p����׸��l��~c}&���N���>��b�	����e���Z7�9;k�I2��$Ѿ�MJ�V�w<K>����u��!N���Fp_�CsQ�0��rW�:h�Sd:�x��~V��҇��7��2}y@�'�B��I�Hg)/�d�f\���B����˔��~�4��iS̲-���,P&z��U��\��]��4���[�5��1�>��d��	�����x%A�Ҡ����҇F��;���ڂ�E��@.�����\I1x�.!$�����VB;��.j�o���-���exZH��t���p�R�i{��>�v�)Bz���bf1�a(�eP�aD�!������gE�4̓�6|��_�K8����(��.6�=��8�(�N���e�����Gx༕he��:���&�j9c��C��:ʐ�V]�+va�[�$� w���'I���#B�7�Sˑ�#���&���ُ��)q�y }{+�XׇW��`��h�׿{��Ś�*5c8��$R*#A��Q/Lǫq������X�q\H��[O��uY!��,�Ef<#��Kؗh�UX�m\��[=4a|�`	Я�\��U���T3�c0���w
?q��WUp�_�Q#��Y�8��H�7�7�ƭN�h�,Ui�I�@F���+�r�n��
4C�/�+s
�=���,�����B���#�����0z�5`�ܷ�Yc���u3c�{"�G�^�U�л�B@�t�u��<��d'5"�Z��;^�w
��p��}5D\T�
�r�22R _��e'E�uT��]D#��i�vA�Xr�$���r-��U=��c��[C�V" <����AOB�H9^���ڂu���g�ۦ���uWݵaP�~��xJ}C�-0�rˀH�ױA��o� 
��`)Mc����`�>�%����7w���](�G>��}t�ٶj�o�H������.��7����u����QI-_�nn���xu^>`��KO2�U~��9;�y��̆cj/�����pswM��2[�P�Hծvyv��-�N2v�/0ܯ�ث,���!^��ʤ������l��J_����_�h������/F�׼khRȫ�WZ�2�8�`��(�d���M\f�����R�.-Аc�7w���]����΀"�7'$���:|,�������]D�X{r�A�:�P\�S(�ZX��iY>S����$(�xr��>�(�?���1er�&h�.��{f;�ܛw�;K2�ԟ��,��]C�J����Q��>�$�M�־i<����(x�f7�����~��<ap7�dl���-�+=�S�Sz��Ŭ�`DerM��ȅ}6ni��V��)�?�`IE�ts�#AD��p0�T�P��+:�^:��7g���dE���о"K��y���K��etYS��<�ĨXb��:-�_{{:�	��~�N��� `?��w֘ݩ��wCF��G<�u�س؁��օ��W�uX�%t#~@	�H'���^��@)@!G�6�z�R(���?.L8�mBaq)ʴ�zU> F�}!9���2� Y��綔�M8����O �N�S�Mk���䬬�/G����LG<���ؐ[��"��z�Z�u��u��^�:������w�*-��j�X�M5SuX�?���1�t�{����~��id�CR!OM����ܤ8��WQ�����v���_��\�1�."y��U�s�$���ҏ�j `��T����N6��K�b�e�@?��o{�<�]N�B��Z����Dc��l6O�[����`xC:YḬ�H��c��I��>��CzHB�e���^�2�G��m~�[p@o!V�Z��ZN����^�J>��^re���	e0(�8+D+~�.�r�V������<ϭqU��d�x���m"|p=�X���}�{����B&�aM)��n�A2]�j;Z���ް{�y�L�n_a~���n�) k�s�z���{T�xw�n9o��W�#7(31m�T����ә �N$�b�V�=	j��ZI=�=��UA#��z$G�4�����_���f�YT�%o���9�%@�1Ĳ���vH�����_�uw(���?y\�"۫z�s���uB���Xm����j�ͿIV-g�M� 40����ж��8g����޻�I��?��ڗ�s�����d�Y^~����I�P������u�	_Q�B���Qu����J���5�F ���F:��T{�R�RX_�	ü_�u_U�P%|݁ed�q����3(�Z����A�P;I�̅���L��u�S}3�`p�2m!Vԥ�jm�׬�7Bm��C�#����_����糐ω_�G���3�I���Ƴ!!0#��p˕������`�@e������j�j!գ1uG��$\�� �v=�r݀S��* �7<�d'`7�̪�^��|�
7-�
�/H:�$��%A%�L������k♥qU�S���g�)E��<�P��&͓����B�z�w�E��d����fC�i�}��:�O�BRX���w�cD��y饍�Y����QIE�bh�2�k�~6��C�>8GNZP[D<wQ�@c'����j��^�u1�Z#*��?�V�A�1�X@�Lz'��'�,͗�n^��*&�>4e1���8���H�ļ���(+#S����v���ũ'7m�=IAD��T4N]5�2�^��*�Ɖw׮���d��#%�e�����ꬩ-)~r���7�:�����8�蓂�%�ن�%6J¯���c:���P3
�^����w w�S���WmׄO�fx�YQ!�aT�[�3����PP���X���ϗ�_�X�x��G+�̶��il5O�2��9�8�f��A��֖	�=���g�_V�*�)���% +RK	�TKb����h6�Qm������L����r`V�TH�ѹ�AW���ޞ�.`���x	uq�$-u�\���� nB(�7&��s��l��2|�VFm�yǖ�����X��Zb�Q���~������2'�@�֞m�c��&��H�V�:=�ҹ���R�0��-�U�م�~{����;9�	�ex7�A
���ݎ��8x�mt�'W8�}<��g�>J�P�i�8kς�y8�ة�<n�jY)��DP	���'|\�)!���J��ҕA�{����^?>:ڷ�H��MD��#f��R6��3�A5�Mꭍ���m��A	Y`�ӕ��ڙHb�>Kҟ-G�r�G۷i�(]�E�q���T�腪@���,J%Z�=�زx������*��a��U�*b8>���o�h����2������{�e��}Q=?�}F���kq���f6ד�!� �cΛ˕,�!Ѿ,ۼ�M��o�9L8yf&�w L���2�������ʶ*ޙ��mh�j��Gr������5_� �υ[�h_N�iI�ϧ?k*�Đ�� \7�5=Hẙc��Q)n,����ݖ��H��pڨ�!���1ziE�%(��A�ȷ
��yG�Ns�r��С�f�Q/uP�φ:W!r��cP�f?�`x�L�^� ��]�4�2�f�9�[��`a~N��EGW�����v��H@�}t�C%�^w̦��i�/���{*�+���V��oC�Hg�]����������~�B��j�%Q�F��wH��Ux���C�C�q5���i�/�&�3[7	���6l7w�,}�.��{�20�M�ʬ5C/�%E��B��b͖��D��؏ ����V0���HX\ͧ�1u�u.�pi��G1�|�����`��k���La����
��R2D�:�E���Tt{m|����`plL΂@j($�g%ӈ�������E��ʢ��nTT�J��^��Zے��0v� �⾏��:d?�ɻX4B�@A\��S-��=�Q	��*�i5�z�;�OgV��~�R�|����w`;\XB��bi�Y��V	lh�:��&�h_���j�Ɖ��ݤu,�lv�s�V��HDD�*��i
:�-2c�N_@������wx�d!�W�#�S��/�0r�_��E`J�Ƭo� �� �/"y��m�V�ɘ^7K8cH�@7ы�}"YԸ$2���!۰dIb�εf` ň z�U���R3Rh&�[}�lq2U65�ڽ_��)�T�2�O������+���V�V��u�>-���)4�J�3�u�i���2�;�+��CWU����Jm�����_eT'Q`�c�^4�|u�:!���}���w���1y_�웄D��1�dvQ6�~����\.��v2��t��q�e��9~���ղ<��V��r��O�I-;�[2	��k)��[BN�z\���e��) ���.5�W�Ӏ��(���4����Βf��K���a��-.í�&ep}�D5�N�#L ��r���5.�p6�<Zs8Bl�t���2Oܞ��x$�ig>�n��Z2�D���U'8���1��QOR�HU>���.�KڴU��w��^Jigc<��� ;R�b
��8!��3E�'���=i�K��B�S��{��O�,;��f����
�D�*�;�'@Г��^�|/���Â���h���k
p�Dg#M(��X��b�Eg]]",i/���D0ճ!ig
�3�A�:�*r��-��d�iԐz�_��l�t�g�C�þ�1������������3�J�4����#D��['�Dn���|�T^�6��}��UÍ��'�C������?N2VC˕�Ƿ������pk�'�{�QC�>Lyn�<->?>*?��������r�3#���3�O�M�<��YYu����qyX���+�Pyr�fX^x���ɮ��H��w��[!K�����Ht+�?��WO]ZL�����6�����/�P��f�%+����}!��L�.�8^�|�:�V*	�M��6:�Oo��sc'��t���x�7�ӗ]��֒.`h���c�s��x`�쮰t��� ������B$��ǣ�������t)�B�bQ�oˇhd�ȱ���Q���\���? e�w��ͱ,�s~��AK`1�H/�*%mt��Jx���M|���ꑿ��;֐�i��C��@�F�#��ٵ���#��>���b�Y[�{#�	�b��I�̬��<��d����fޕ>��0����Y����>�cI,`e���̂NZT��_�#)�L�j���������Ҟ�����e�M4}PA�m���>TQ�?���耢��I(*`�]��E�"kNҟG^��0 6l�i��{���)`~v(dK��:��e�r���B�.���zP�y�We	���Cw7�0�e[����8�a�h��ڙQ���tW��M
Y�bd��0�q^'!o��Iz�����r:��8<�V`��}=.)���w��[X�p��#gr�N�����_�4O��BPp��YF�h_��h�Y�K�&�e��gn�-�ƺ�����V�E�Z���I�Jh���������#Pݡ�J�W���(3+�\"7J��X���\�Pli �4k�;&���l��p�R��YU��>^� �*�� "F�Nn1��z3�.`�FY�)�7s�u�j�_�-4��g�����S6�T�x���p3�j���@'_0�+���c=gcE��(����A+���W�����.�%*���bs���{R9��rs�R�E�"���8�Q|*���<�Y̜��n�S���������ϙ��������ZF������Q�����5B���=G���ڋfs��W�D��7m���E����$����]*�zmfW+C{���D�x�o'7���y�4��Zw\Z�Y�S<�E��Ap�#��^�u9���޾�K�	�C��V���*���[��/i��p�֋���P:�U�6�v��K53ե��Sue.�x�v#�^rԜ�U,���H_>������ڣ��H����w��{�A"�v�3�S��ifx"Z�ﹽ�:����9 �ҙ�l)/�Q�Xo��f��� ��/U_��r�OG������t��~7PB���"�y?�k���8�k�]b��qQ}�]�rLH�\�� lϙ���Ӡ�e�'���iVB��"�孵��z��9,(JR�)]V���탘��r�g��$^2oy�u��j�|iV#�1�5qF���Jt�ݯŲhWXe(�co�[���*��i�n#�ggϧ��=�q� � �;�N9U�<�.j�������Ɓ�mMZ�B����I����m�ZZ�r���pR-�����dW��@X����"8���x�}��E6Za`�H�炼�h�cL���o��a�y�G��'��}��CaIX�vs��3���.���������0N�-9!�p�G�Ç�fm9���z!�q�����^�@[>��N��v�avO��L�x��z�8zXQ�k��:�
\d�~�`XB�ԟH���k*`w`ݫ��PK��&�2x����2X��>�(�~���%Y���.Tz��5���Ag����e���p"���B�~y��Y�4l��4���̪����q^t$���4>`�&g��o#y���=.Wz
E8�<]�c��	D=u`���7�H���%�^4����gbՂ�Z����r7l��8��־�Q���_�-c��l���ǋ���-�?P�����{�^#�:����!/����-�P��J1���״��X)�a8�n�X�x��Z�� Rnޘ����E֠B��j��+�ET�y��P�y�������̿`[}C�潣����j�b@�����Z�giF��Z�R�%} J� o�/6�R� 
�Wԟ������gʄ����#"��8U����@�WA��3��p&3�A���@�+Jl��~d����\��k�HS�&�lT"��7�g���a��۲PY�\�n�Y�d9\��ܡOc@@7}N���MH��z��\
اݠo��dC���$r��I���\�5�������D�= IY�ڵ.�f�����\�����ag�P����<��Jj"��2x�s�e���"���`񨙌)f1�L��_���i�hY�:�o[�;�q#��P��rqK�N�>�'Q!�C��!�����fny7_�,�cl��x�V���#3�2���A
�Q1�
�=V��q �M��?tU��[&���4�h�H��C���gtu����H�KJ�w��2�4P٣������c��'�p��Ċl�y��Ma>-��l���V#����b9.�R�o9Nr'HU�̍�)���># Dk��8�x�$�Pў����iRH�r���~=d�^DoƩR	��.�*�`C��A�6Z�^'�� 
������j�r�0XV�W�I%c�3�L Ǽ_���i�|��/�1}E��v�B��M9T�
�=:Gv���$U�拗���c;�'Z��g
]�k��|?��8���sV�k�ɬ��,���j@�ԦU����~��M��|�_��$.���� ��)���+`-TQ��~Q]jFE�/o�ԩ�1��\��_F��[Ԥ�z�W�U;>�?̷���Y�����
����_�za��J�iG�|F&��F��/�b�|rv?i%�)�j���#�Zf���5��gE��ȹ�_��QreD�^��	포V��J��.�����>e%�Z�i��)�}jܧng��>U	��՘&
�����A ?X����=	�=�J���o���"q���%�s���&��}S��W�/Jf��o������
�<���4�́ۤ�-�>'�D�ٴ T������B��o��m��Z�8v-��TG=+^�sJGƣ��qC������#�/ܿ5���Ʀꊒn#�F�-T�(�V�����p����,���Pc*a{�_��ȱG4�쥜5YH0���8<u��+�[�_���5�Z��+ov�=����ff�u��zz��@��5G��������Nqz��=������!6��ox��]�[	};/�1��ق�ϛ�a�����^&
�ML�,�
hM�G'D͗n�W��Z�2�jZxb��g�n�B���l"K�0�`� =��;cTHgN����ޥw�%z��܎��\]~w�����*�m��%j'�,dV_mz���g2�$ I��`���n��TӖ��KT���7@d����_<� #1h��<?N���
�:rq}�)�n��s�.OO4�
�[��avݔP8vI6e���=2)�U'�ӣTZ��6?H�l�e_��BqŲ���ۥ��RqRP���f�����r�c �Ɠ]yE�*�����ȀY���	�@$���]�%O��HN�l��9i���}a����$����n]g�ҷ
��ި⩕C`�7�B>�i�0�%��/S����<@bm�"Phk솛 �т0��MQ{*���Әc�5{�J�4;9-*,��w��j���΢��M��뎶$dS�m�鄞�.ֲ05���^ԁ��F�Jn/d�罄(��cl����U�@$������P�_cY@NJ���l���kB�L,�A�Z���ͧj�"���]��A~��Jd������O=���]�t}L�c���`�4:u#Q��xqd��XXA��E���E�����V���҇��"�ά�}�t��/�9Q�z�������ZvR�G0��֟��/M�d�掺��]����yC)<�'��HQ�..���ɽ�N��Bi5�@W`��ѾV�4p�2��{5U?�:�Ѹ]v�1�m��rR��G8	e�Y ��+s�}��" O��7��&��^UVX@�j-<��j�k�=�َ��j���'2l,�o��I.B��\VVüe 6 �ݿ�-��<�֛���<�<p׮b @ĺ�n��6�p<�&�N��I���E�P�<Bhm/jH*���y�����+�L 'һ�����#�b0β�)�ᨏ��:����Tݦ�TZ��ii_(�ϊVS/L1�p�K�	d}<�XJ9Vk݀-q�W�D�jn�}�'��aH����O���G�j�������l�;��A��%����ɨ����/uQReU���F�\$' ��M�s�z�G�Mu�n�u;.�#f��̱�W4ssI��������s`���vY�'�@v�g�i�:
tR_q�RX����µP����C�QX���-�٥�qF�rd%˴pq���P|�����\n�c��6��.�q���	u5}(q��n	��J�go_�(&K�T�<9`h�\���CI6�Fei��ۦ�Ӯ+�$�)�1:s��$�\�y�2B���&�ɹde8�έ�̭�w8��%�Y-�V���yK�����(��{�ެmܞ׬,��>m֧�vF�� �p�-��B�tF�)����o���d� S'�>,��ul\�������v;��w"�e`u�[�vv'aA�oŝuk)��~����0k�K�����b(�U�lU5Eک��'��G��?�����ZX��=˦7Ѐ}��n:tN�nso`{�Pr�l��B�1��{�	�e�K\"�u��x��譯���H�7\���Ѧ.'�k%l9���l��`Ֆ��Qɭn�Ǌ�KX^Cן�ͫ��9��~�O��,/v�7L�#�^��۝sf��wk������F� �y��+����Vؘ���n�n�=.H�I��C��f�ڂ�`�Mj,P���#~����\��x��}.yKs��R����<�
 ��U]	�s5)3�	�
w
ffj
n�>��ڥ*�5J�VZ�1K�L�j'u�@s�C�9	@��r��5�[=����=���dz�ڪ�hҢb�T�ˊ��f�������	ӯ��Ë2�]x�8�@gu����CA�1�Q}=�t3ARb=���y�z����m|F�}�����gS5E
-4f7���a f�XnG�jn!�+�`y���
�E<:��7���JQ�����Lp���ε�7��J*{�a�4�Ԃ����6g.8�f����/�������{yC3k�'���� �o�L�kH���0찀I��G�x��"�&������[YDL�
��2\I�|�H��N������\��4��_�)�m��x:~*�Q�K�΍,8�u�b��s�4��r���:�{���yz
��`ݕ�Z
)8^=�zSm:E���aD6ac�n���Jk&Ǐt7|��D���7a	 H b�X�I�tkw�.��a5�<��[$���k�S�
�D^��dȚw��~��ꦄ$�6wZ��)it�Z���y��Ph`E�^���`����#�B`-DkRIy)�%5�]�P��=���-a0MH�S�Qr�(���Bx-Y�a�_]&��V���hQ�� 0ET)*�I3O�n\-��;~O9�<��U7ݧk|�����gy�٤lzo�V�I[TD�@�K�'ň?s�cJc|w^h�_�-`�����9Q�Vb}��G#=����v� ���R�\��ؒ�Ǭ�:�#I	Q�S:���[r�4Ļc�D���ŸI����"c��E�䁔�P��+�Jß<x�|�p��@h��R�d���0i� ~�2��7W@_���=I&�<X��RfrM�o����-lG3��9���]�q ��P'ĳ�aC��2|pv \�.(e�zF�!���������P̕I8j�mԑ�U��T�xǫq����*C<_m�N���~����q��� �b�h������jK�1�]��ح��e^�E��:�/�5� E4 �Z#�[-��.F(y��$\���.�`8�f�c�|.��)%.g�k1�ӕ�u;�P)��E(���=��Z�����▮�6��t@���<���E4���Vmk*B���)ڜ����y� .eq�!���P��Gת������J�M��U��ԉ�T1�gbW#Y�aw�����:)�W
>�A»�%��!��R~�+�@q���ۑ絡��F"@�zǣ��
}�LU�̠B�)��S����z>�J�C�ezIE�Xn����#�~_|��߳���?�H���J]A���h���>�vT{fT!�(�Rw�Q�p ��'�P�Q �4΂)o%~la��$b��8�0��XiTi����i�����h?��#��~�X)+M	����p�d����Rʡ7o��>�V�mؚ����{Y���'�� F�u&#�_��=P�5���G��O��b��x�>��BC�)�o�,͕��i� ��Rz�Z�Iu����,5��F�_;b�2�T+:0p�����XH��"��m�𦟻G�0^���]�z�f�R��0U�h�Q�w�oSp3E��Å���R���3|�!�O2��"�5LP�C%L ��y�j���)]��o��.t]Ԍ ����4Liw����le�ek�Pq�b����|�m�<�䜓��]f[�Ub��C8'w���K��,=�}2EK���b�)v�h�ϔ?�bE
*2��0q��w4}߉It�c۾��:��/L�y� x�1L8^}�|��} � {&��['T.�b(�|�	!�7.w��9)���>�g�����rR�����,�h�îa��{yt���8KxNu
#�/;Lp��׋�yΓ��!��ٔHz�d�k�
u>���s7�*���곰���HY�V�� �����T�wK��EH^�˙ǈ<<�Ӹ��U�����W��_5�b_v+E���|c7�����4�L�k>�=�@�6Hwy��Q�d����n��A�U�8*���>�[v{�L��r�A�ꈏ��F{�Ҿ���3E�x"�����v u0���={}��b�,�Np�P~�54�_	ұ�����$؇��	�qz=dw��M���9-; �K�>�}:�ҳ�����M�x�-�률����p��.�rG{�jB�U���PG� ��V��]�-��q�\��Cf�ɫ�\g�m��f{� =5�_U�x�3R���]�NL����)�4�d4�Z�ګ�#�y��cmQ\6�+�׸QHi�!y@��8���2e�P5ܯ+�e�#��|a�����z�>�t�d����*p�p!��m�}��zE�  ��2�R)O�o�7lÙ7��Px~;��cf'�/E��f���
kn����v�|A���ZD���E��ly���1�FI]�M�N��b'���Y���{���h�����~�������H?2.�E�:���|���^F%^y�V9��[�"!'Ejwؠkl���UBؒ���$K�ob�\���r���:}�1���=�~�J���2�wat��r��e5p
�ku�nUu܂�4�bjoO�sʍ�$pr�|!��Fz��n�&�KφIp��Eo*(�Mf_N&��̗��,�B��L��5���R�2�����~+�`H�>R�w�qm�l�?6�7��|Z(po|�+y�]��z��®d�	J�8�c�h�/ť�Տ��>V\BG?�1_�����Rq(�躈	�J2�?��}�z$��
��O䨿��)4s	e�;���wK��)ie0��U
8R������NE쭙�z���?���	3�P<f�0���R���q<�x �G��<U�s�����"�+���(�u%T��)ȽW)�<�Ǽd�w�[5�@�\�e�|�;�}�������w��[��������� @���D����!�����q�Kp6x���'H�)ޅ|���2so�L�����d���|��d������q�1�@9��!T�;7�mm��K�2e�a��jљl��g�ĎvU��cE-�k��y|��E�4bp�q��+#�l�߻q~�w�9��F���xc�/�Vh
u;��.5��:���6RJ��h�R���������o�`qĆh��1��z�8�3�rN��@�^��-L�W �J�6$�)��D�6���Nɕ�H����$.��2�Q
���0)��b~�'`�r��QQlһeȾ���d�ԏ�}�K:^[�\��`/��=�q��#��9�����W5��!���,�q��� 2�iJ\KS�<�݊�@r�Q­���H��ڹ9���0+���N�9ⶫ�	�ZGg�T.;oW=���U�eK�gS��g����>��B7��%k��'�T����9� a�L�&� 8�A�@� 
�	���Pv�Ja��|�~d��H֏�e7�	v!|�k�CL ^R�4�V������Q�X`�6f=��&)L�Zx��ż�2�z���2aS�����)r�3(�S��X�5���i���xF����ƃ��IOֿuZG���S��H���w�k�%�#\�"=v�rk�� ��1A�l��|�.�_<?��Q�%�0$�S|īS�	��=Z���ϛ ��6ٜ9V��`IyG�����!Y���0�L���0q��K�][�X����:9zL��Th��&���j�c�w�]!#t,���:��i{�E2`4��� �[��]�?�3�)��z�3k�G���䏷ghXw�~�E�o���+�J�W���EQ]}b�'�/nE�B�g����agc9�y}��~>�/۝L3v�U�'��{�i&BX��zH�2�!Z%-|EC̞��������r�:F��JT+�U�o����=#�_��_u�(O"\���yo�C}����&��9��@a��y0S"����(�OcI"�_p�"���#�}$��Hv?�/��=��8�g��OZ[�[\�V��f�G}������#P��
^��s.�K�V�;���}��L%:�z�����}��h���� ��Ȍ�H��!��f�嚫u�b��k�?���VH�w����n��h'�AF54���֡im�O����~���D� lPy�e:9�>�Aq�>*Z��m�,<��F=��u x�TE����nN�I^���w�EV���M�����q��t��V)#]2{(Ƅ���e�ˉ�)��y��f%��>ڲ�X�SVm� ߤ�Ztq�k�24k��<?����Ѷ����jJ�X��h}�⾠��v\�STaq{D�߮7}d�xfZ��'C�9J5V;���Co~���{�S�d5�N��h���T��5�@#欷W"w7^�C%l�*���X��*�&��nsu�~��&���i�w�0�I���h�L����`�Y%i�>����81"�J��[���o�{0�Qa�a	@��"�2��s82��5����/��^�<�FU����h�h�́|�yWJ�Ȭ]Y�ŕL��U.�מ��D��L�C�oZ�B3�&�J��eDD�8bm�����8�X83����ǂU]l]n��<� ����)���M��gI0���xcĹ.����L��Ը)70��D�<zs0�R�b�E:,�qF�r������(�6a�U��@�����kV# M?�%�آ�t���A�*�:�ac)�n�� ��7~�N�F�j>$���`����Bg���jFk+���OO!J_��$�Il �����ٮM."�o{��H�5�@U�چ�iC�Q ��gvǼ�?�`C ����+8m�o[h_�f�]±:�OB�Kt��5C��V!oi��M_MC@\)��j�?n���I}D��m���/��t�M����p:u�5���?k~�28oK� ,d������`t��`^����C�\#
]�7a���c��/�:� s�'��xw���\ί�`���DD'�$����\`W�)���T*?����/�C̿��E6n�;`�J�^��:ͳYzL��nF!���T��r7k(x	��k@��OueE-*d���N�戬�5�|�j>�`�	��]��))����?��Xyh�ȫJ��@�&��p���j�Hao67˟ E&��XB�vE�852��M�s
�GokM5�vx�^�5}1h	%�0&�ݨ�T���:��	��62�kt�9���B�w�A���BI �4�U�Fj�b�V}fS(�}x�#��K?t����3�y�K-�nr��7VC[�V��}��JD��lp�����9R��s��4���;
�U�G%š�>T�Xa���2��ޱ�mD�{kɞ;�y0*|)�����7k���N>e��s8��!y�k�����'�j�۩�Xa���Io묰�lN��\�S��9\��o�f��F���M���t݋��4��W'c�*Ԗ�J�E\A���!C\g���풨�(�.�^�o'e��'�)����wإ!���޷�1��t��.�\�֪&:�`��� <A-��$����ؽ��a�g������=F`^�}�ey��h��A��.�|ыǨC\��,K��ڇ�KAE��a�l|�����F�Gv��E)��@�8N�\�$9H͑��~���!���9�����$زn�� 5[���#�1q-�׬�J��YՔ�2��IPI�IN#ۣp��U���Zg�Z��V%�tPO����	S��B赖q�\F�Z��[���(�v��5W�s������A����s�4@�tiE*����a�F@6.S�b�w\^F�GN�t[i�B$��-�:���A��������B�X����`��Tg�'1��[_��u��(�5;~�5��⧕W�v���;Z��u�"L:����A&8�7)�|�wXƁ���\�����
���7f�p|i��oM>#�!/�`d��0�%8�7�Y�)�9��{ə��)������R0���}��yYħKBu�Մ\5����e-:�mTR�&@<&&�����W�|�"��t���Sm����C{T�z��{lpL���h ᕑ�-����ykxPo��ݦ��$JAR���Dt�ޛ4��l��i��'m�'@*K�dR���WH����JU[�^�ʦ�b�	�1|�Rx�wX�U9�I׃vۊ��B��~m?�$J��M��Y]��v��l�r����4O���lb�v>���4����z���A4��#����f��8{����]h���0]0������r{r 8V{�_��o��m����9�$���h��&ue䞋V%�;g��̘F��"9�8�/z���c�;gXX#�i�,�����{� us�0Z&�g��}w�ֈ��{��+��/�ۮ����̈́Kk,�j
ϑ��Ѵo;L�Hh� ���4�}m�j�o�at����"��<�-�t_�����r���@7�pvU���
�0����$x`�vyМKȗ�Y6�UH�0�{Y3�𦋨��ţ|֦K6E'yLU��nN�-·\̌���n�\�Y��\N���{]}G�a?9��{���\A��Y5�A�%�����o�+M!1I���JC�^-�'�"�9WY�}��N(���Q��"?8�*�)�k��G
��6l��"�َ+�4� Ȋ�6���/Y@;��lT�O]&�S� -d�׺b�{O/���N�'m"5e�	��ԭs5�j�s�K��@�a�X�
�O~����!,6��<�m��~�F���\HF���ht�n ���������)Z�-U�{:���1@�FY��ߥ�Yx�&fJ���W�ǡ��������!K�{Ѽ�ߚ#���v5�{�(�W�د�J 5���h���`��^�h!\S�����dF*�/��(5��c�\1����к��"ȫ��r2�ᅗ���{)�晵*!����+�.��J������rP�s"�^?,&o��f�d�$�.��s��5+���5�h��M�F��<��O^�o�&�u�+!s�쨁Q�s v�*x��e��E��Ƹ�$TӜvR�&0vC8g�E�T $n$��� ���UfǊóԸ���Bb�VT��u�Œ�bU���1��	>d�C/��"5� �q��~)��#2ì?�.��|\:�ZE�q���V�8��X�I�Câږ��Cs�E"�,k���~c�I�������`��94�Ww7�q�eS�l-۫G�~&0�AbJ����sMR3�ƿ�A��
�$J?  �>wm�<L����sB2 	�
���c�Ȩ�J�[�?��֎',��y*���7D;���4�u�ɴ��F�dy�e���pk��5��Ԝ+8ߍǋ7sX�v��o���V��ͭ�61����W�����E�8��\8ޘ�7��{�4��KD��<d~��*'I�=�w@:C�5�MC�E��<���yׂx�+x����M)��'Vz�I(ݠx����A��aF'�g��ܑ><衖�����wQIx+$Ϙ���5qI��B�p�PI���5kA�Ԏ�9~|��I�X������?���������˚�%d�E8r����ٝ:��Vq(Ȃ:�'��aWUd��~%F�8�q��|MH`{�F9L�m6��#�z�u��΋H��X�?�j#��B؄r�Kq���>P>�Bӯߵ%V�gz�����M|�e[�.�_u�:�a�pᖬ����W��V1���]�f�U�1%Sb�S��R�:� 0�V��3}*K���1�]�	���&KX�:�5ZO6SV8j��+x҇�z� �]}�~)ƕ�X��~�^к����<��n&���Y��+q�LՑ��V�dLq%@ɱJQ�1@���F�'���7������?v�U?�Y���k
��ck�_�a���
����"eW����R}aSc��O���4���!&?n����%�pj�i]������#<�.+;#L�.�_��w�tr��E���
"!��v�9�Sq�U7�y��U��Y x�V�}s��ܪ<��a!�S�?��!��H��cvׄ6>a��U�W�3N���؈�պ��_�ޯ���=崨ѐY� ����'��t�%̊�(�_V��! �aX5҈U?��}9䁊<�{�\m�<�����LY��K��� D2 ���I����儙�K����6�w�> D���I��bZ���6a�n}hY��f�}BMg��f�[�z���Yʁ"�p[z�+����C�1�]I�8�ۿ���s~&AX���bK�%��`�uu]���AV�F&F��eݡ3.<�4��3��:���Da�y��I���\xeY�� �����L��+V��{=���j��'갛�f_��uK�x�B��3d\�^�cǖ*vL����b�i
|%��!.��;�ڕy$e���QHi���>�ϓ�l�����炅�8��{T���H%�����G���K�!���V�W���:�2��]cTHW6���Cs!e,9L��-;�e��ՍWV<bR>}�?�|:N��)R�"���KC�t5��m��zL�%ԋ�h�|Wj�#S��fr1��u,����bK��p�In�V[�L힫��M�Z��?>�c���M8�בܨ,���>ݻg��������&�P�f���6�r�#j�'�Z�UՌs���6�*I�"��g`���Έ�&ژ�@�,(�ֻ�Y����F�6L�>x"�1����7�ni7q�v��G�qO�����I�'�uw�f1i�ѿ��i�]�UiY�.Jt�5��z��(�����!/��Q�%��K��N炰@bqo���L �0���fX���a�0з���������gWN�k�u4z����,{|xz�Pl"�%����Dd��Z��ҷ�k�! Eu��5 �Ieϣ�Xu0��Z���M�W�S<��@�&�Y�%"<�e&�}XMyQ�#��=�ϏS�m��g;����fr:��E�����3g�۬��.�ψ�9᫳�!�A,��)��7.����QE\;�&���{%������7V�!����a�i2}Į�4��@�n����2)�����9�)�����Z���7J P���������<:�J]�yt2�e"��`�Lt��Ah6S�R�\���y��{C��������$)M�v�v��vE�+	��ܴt=]��˘��ʇ!��ˏ3������/z���1D�T^[��o.�Qy�Х|������"+]2Z�Bh�����yV>�I�:�-�hs�]x�֣��[M8-0T����:N�u1���G?䮶%��I��"G-��67��|am�>:.ʀ���X�q�s�yP�B3La|���9�8}W��Ǩ�7�X^Bě&>�!^��%e����;=L[C(�O?�mZ���p��@rC�ʉN~z�H���K����#9���9�-߁��s�k���kd�B����# �`֬��L���:0��IG���hB�m�O�I������Y���B��#A���h{W���6�j�3���QpW	u2�WQmy��1�u"""�m�z����L%���b�iƞ��S�c��_�4]��qUVW\f��@�I�{��p�uS�$�'�=��:ɱ"��!>A���G�3���4$h�~sX�*M���s�P���8����;q��%n	D�QT`��+�J��ؙc��H[J�D��+>�E7X�MBNE�	
}����D cy����l�
�E�"�Զ�D�&_B�!9�0T$�<��$�2��̖������u�g�"E�Tp�O��s�?w�����e%��d���9����4��OK��.���}�E��Et�L`MQ�$��?Ȅ�I	��)���r�=+�>#����6�]��=�ţIRz41!!�]з(��x��]e��Z���/�������e`ەT��N����B(��B��/��m��5���Tnk�j1NO>��thX[�q~�*_�:y���f}��eP
���gL�b@�@�m<RfÔ��o�)HK(�&Tt|<"H+����yy�׾�r�ɉ<~��d]�7X�(J]O����GT�VA��Z2��s����w"���R,^-G��Z�4f�`�l��V�} �W/B���o8��R��Ub��i�������Ԉ���D
���s�n�� ��i�X:�4����>�١��o��4�r֖e������hw@���"���uK®c�_`Ü�0CJc�A晜ⅽn��:�1��X�"����^7[la!����m�a�*$^^'���*��¯n��;N��lԹȔ��������SB����ߙ����Ņ�UR��-}���<�C��K&���u�IX<�[�uF�F��a�w���{lO��E�,@�9���-��Y��K�#�S��~y�C�\��1�#����́����|I'�ۖ;��İ�U"8:�]G1��j޹V��L{�.Ka�	�l������dF��+:8�a�r�>��dS��-a�G4�kZ\�O��ן:���ƛxڛ�S��2ʘ7�˞�������>/+pM7�	A�,�xem�.	�5��l"�eWQ�q�Psx���=F:hH���@#�s)pB]�JS�.7�b�C���c��]qF����g�S0��5�G�̮U�؜��a��U&�f�OB&	� ��I�0j]�2r �&3�s,�����ԯ�`�2�w���m,F; >��3��R#���]J0�HE4� �b�f�r.��ꯂ�K�2��'TSԊt:�^|���{�3��Z1�*8�P�9�Jv�!z$�֕��u�M���o�8��|�y}�ym'�k������ ̢��zU	�Hs�z�4�Y�K� ��NSDW���m��yw[A����3$���,�b��L��"�3׾*/V=_�%�IW��Ѳ�I����k��o}�f6K����>��=�3*p���U��+ɭ��OY`�k��������B&/,#w�b�,HL�ӻ����´yx�5��9I��2[��ީ�	~�V.h�;��vw�<{�Y���]Ĳ���W<}�X��/F#�'JCf��}��FY�Ƈ���Q,�*�Ц���C �p�SfM~��,�S�\�X�8��~�_o�fʥz󽹖S{���jpŦ��)�*�n��,Z$���߂�9*Ű��%��,�5��&6��������
��ݗ�6'�m���|.�:���ï�ME�s���0��5�Es��񘗀���	�5����gc�C0���}�;pF�R�^i.S�f$������Z~e�n��Nb��vL�M��E����e����/��B��y|^NK����Du��F��>g.��$!IWI��n�����1A�i�=����j��OQ��x���[N��qSK�:���E�Q�%�!��k���Zz�S5�:�t�;	���׳@�e�X�a��5�e�)v��;2���F�:0���#��!t�[ �O` ���;�4�h��ֱ�:d�a�����5Iѫ�������L�����g�\
�(=S��Z��*�K�QJ����!�	�M~��TӘ���������p���i8/�� �4q�)j[W^HB��.�h��܃CT�ፔ
.e��J,�.��)v0��c�i�P�fق�ȣT�� ����������5C�%ܰ�ʯ�r5�^xST����ߏdhT�&�w�`���S�s5���x�T�m�z�yʐ@�+o-��MpV[�����L���!�����#��5�P���q8`��;]���Q�:)4tT�A�lN�v�*�=?`��B�_�Ð��yk��-/l�4�ַ����a�kv�}\�T���>�U��i�ʦ�3Y��L��߁P�X�8��o��ղ�j��󌵵Kqhx*���Q��5�Ai���	 A4������:w(�\���bM=IOm�Qޥ�)��+ì|�$ɮ'�]&��AFL����f�W9�N^�	�.�#G�NGW��1�cD,��P�Y˳�=si0}tS?���,��Tm�*h0�qV"��D�X�wQ�<��PDꀔخG���l��:JY=W}�TR�n���v[�4y/u���]��*��u�G�y�by�bq��"�:���w�A
������R2D��*��,<�	�?[�̢��h����c�r�(�Ά� *��"��7�ܰ����^�����`�oխ{۷�фn�)Z�л�UB�N�+/���8� ��چzs��w�>�5q�5d_I_��������/��f����n���2���������%<웸l
!�b��t]����+$��B�d�4��v1.�@ћ� h�p�6�2� �~9�Z|`��\^LZS/��C�#���-��F�d!�R��W����ϕ�}��0�枴�s��m�m�L=-������z�h�j4�>&j�
�����`��5�ޅ@�%U\���8&m���#b'wy�<���_�R:K*�G]
�$���Ɵ�˫���ԅ��a�H���@��-�Ȓ�X��H/Wڧ�ڢ1Z��/����vK���B�ʹ��T>�{�3ZO��DD �FNǬh15╀���G	�-����hZ5�����$X��#���G3W$;�rT�0���ͭ?:G���y /ت��2K݉��1�%6鎂y�W�5 W�M�H���?�.y�4�"ѵf�i+?.���bƿBb"Lͩ}���3O��`��z-�m�}y��C�$q%�俉�&pR�+�j�]�����_.s��PKǂ-�[}X?���D��k#>7�Y�:����
̷V*�"v^�j0tPs�&J�U���e����!�c^��9�}�<{����I���U9 @��v�������&b+�����y��z��y�	��~>x/�a���g�l/S�Hf2;a�ʸ����Ŏα�Ш��	�R��7?$�D ��������j�픇�y��D��"�`W�j1L�?~Fn �������F8�-����m��kf�\b�AW�	��9G�S��>�bָ�M�4�;N�U��P�� j����?�܋���o�w�a��f�Ӱ��4 ?w ^�U��-V˱@�?��c;��F�$X�w�T�:@D]�B��6l1\��(8�l��ԹԠIm������I�56)�h�<K�����Q�򘻍�����/4�v@}��G&d.����ش�j"{��rߙ��e:��|�&��zBG�h������$\�~�HT$F}��a��T-�`�6)�A�e������N��R��;FUIǽ��h��UB��g0��ퟬ���o�n�r!��L�����_>�?y�Տ�3��Ռ�XJUށ3=�p�C��h�ߑ�@bNL%�5�����>�oT�r8p�s޲���E-	,�D���q#�r�%ޱ�61�<xQ7�N�w=�ʑ	Ed�-��Q�� ~�JY%��5�+���麖p�1�QW��MP4�'1�~Ec傯��ԃ�Nt���.��N��y/�Z2})�b;6��q�I�@P�8�����QOQ�>�}<��Ү�z
 �KPtz��$h�k�Rȓ���h�ʯ����Z���${\���uBH���'jG��Gօ�5O8���5/y8�}B3���/v�_��<�&'�O��=�f���HV���	ORk�4�ӂ���Bb���Vb	��7^�|�?��>�1E����o��O��qg��Dwj$z�T�А2�lL��L�B�qwH�X�pu���A4��Ԙ�l$����ha��,��d6[�"?�+�ibl���`{/C���`]���ۡ.�о��ԜX������H��0�'8�?`ѹ� emђ5Rfk%O=D�e3� �V��3���T}B!�;�ZW�E<�F�.��ق��$GH�S<(C�� ]1|!��\�s�b�Qk��mL��:Iy���?��+z�G}����|E_^�޻��L��Zq���g���x�h�5 �`X�w&��r�cB��Ů�Ӕ��+���
s�����\Ho2aXA""������;x]�R������{=��l.U���<�����/y)q��s\��" ���h�ݎh����$�r��*h����6�̻6��{��	�2�w���~Ȫ�͚G �v3
�mV6�^�����D�p;Y������V��!�N��~�UUtڬv+��p�Ϭ�������U!@xCNղ����yIS��<n�`?����O������q�E9��nB!�d�esć����.�0��F��X�Sz0��!?Z�������s������fp��&��ߓ�U�qpQMۍ� �#�[�,�Α����8��b��tk�V�طI��x�9��i��Z"��w��Gz<t	)>ry��t��=�a'D�٧��4�b�Ӧ�}B���'!\ �s�j�nS&k��4*����FoO � �71Lm�@��_���8�9�B<��$QC�����:�E9&j%���n���J%�m1_�}�*�D<7��笽�{�,�4x�Ae��p�L�|�iH(�H>��U&�V���W=ۚ���H���e�b�l9o ם�gT�|�=Z����tX�5Ё%����'9�M�*�tK*k�Q�Z���p�����!�9�,L��[ԛg~Q£鉇Ů���>�rk'_��%��(?�\���z��z<W��;�A��x��K�Y�v�9M���$��&�;9����g}��n&?�4�-����C0�	����]A�N*�:�ǣ���8O���ψ��p�U�*��v����ii���	*�ؔ���&Sr��i��%�r�Qq�M�Kej���5'"��Ɓ�$^�5X��Q�C��xI*��ڑ�k۪��+b�F@���l���Ј����-9�JO����K
u�(���?�X��%�b����4FM�J�I{���0+��i�5N(D�gY�\	:Y>�1�.9̜V"$t|�����s<��Q>�v��7��	f��^��#g���)Q��{V�/�0��>�q��f��ܱ>&L��|n���vd�Q3�����,.d���S���`'�,Wӯq�yv����������S����1 ��Q�R��Z�u~��v&��&����:��L7�%�\R���}����b�Ɠ��'B�Wq*zsuv�/Ed+���eK	G8�v�4�:��Ԩ3��g�t�c��������a����bD1�n�t@U�h���OĒ�ͫf��>��_�p�?��!
�_���q����=���x��
ʑ�M� �	W/�@�kf�2�k�^�/��ȑ�1$2�\��옙�,�.��w�w|J+�YK92� �I����K�B�\㸥�n���%����)B�2B�/Ә�F[A� �rյx���TA��Q����ޅ�_�{�칷��u�ȵ��=��c��L����I��B���|4������7���d�v�����^��������(�SO)L9�</H��^l,�����K��?F�T�*d]�f�و��lWɪ9:?�B�]Z��p�ڮM��/qf[�zQ2��|/26���#�,�HBi��e�¢�v�(
R 8g�^�i��G���Cv	{�]�۳^V�FM��x��*�4p*�oN��$Y͡�#KRU����rN�KG{��o�4ꔢ�C���m�elbv�a��d�>�^�V�>0g�2�*�C�9�O8��=^�����S(s��Rl���hc-��p�7�E�te��Q�TPY9�hN��=apv�6a^~&W�T��q/9�;Ջ�e�jWmX%eiL����q�{di^,�?-C��
���/��@���!i�n�IJ�)wpG����BGc�<�Y�ȼ���`E�˵�g$Ԧ�9zP�\� t���U>�HW]�̈́�{`�H��?E����֯��~ٚ�oAu���@M׫�s��
�yl^gf�О���9(K܌P �i"��R]3���U�T�c?�,��$pe�!�$�ܷ̤�&��̳���f��O����ܽ���Z��L3�)Ȳ��QA����"��O��<��?�}̈́�t�{],L�j���2�������e�{����D��=}�Á����	���4*53r�<�n6vpdy�*:�5��F]I�oB�,���0����U�Dڀ�x�Z���V�l���~��͖��	(F�8}9f�.;VUc4��D�Z��Y���{ �f��l�c֤m]��jy����OK��ç���d<�&iKE�Mϝ�@|�y���x!o�{V��<ZI�i�3|G���9}00�v��w�&{T�p'&��Ԭ��Ab����đDB��0�0�kY������|4Vh�Qz3ײ�=�ի�N�q8�+96-�|��֬��������鯷?Wx�~�W��H�`˃Z,�����Nʊ5�=Z��\@E����8 �-4��+����g(�ÖS%� �4 #݈�x灋���;��g֎��j+��>�6٘�>AFrLh��[1o
P����W�6w3&g Q��Ο�����{���]'X��+V���#\�8I'��1�Oo��A�-z�S*z��1�8�Z��Չ�V�e(�j��HK)]/���7��o��9��x�o�I$�����)�&���K��ǀ楳G+�K����q��o��։���t����W�X��7���J�_��A̸�i��є�)[����O�"T&�֢#��'oǗTB�ه3�YtUF�B_��.9���"��C�8-�r���
�(�x͋�_(v���\3�5��$'����xz���>��5����Nlf�0�]�	J�����f�sx�a$ ѐ��������W�c��,�y�*�����4!�8j��`�U����∥�����,��Y��}W�!��(�*��������l�����ߒ�R�Y;�{�]!��xPF�^d�b���� ��(����PE��>�+�Yd	a���n]9�$�w�(F~j� ���x��q�Z�1U>0u�B���q�W�2ŭ����<��2yQ �g����8tdY��Dl��P�>�aV4% 5�;��3��S�	y������T�[�_�ŻSI�
-���WÉ/-ʘ�/K��3���X���,+Hu�\�ӥ�8D�¡���O,#�AK�� ��k`~Re=~Xc�q����k����t��TB�>��5��X�SC(�<��Y�!��2�Fe}3�L�� !M�V�9��~'J/��?HE�H$F��9ϕ��+�I�(MyC�s��9��3�b�wz�,6cr���%�>��^�t}MGh�-�8��{M��l\F��t�6�з�à��z�l����$��īs�b���$,B6�� �AXJ�>��pR�:?�G�+b��ߡܹ�5���uZ��/���Ǖ��б���X�U�12D��šY�����(�1:��l ˺�Ԥ�3��ʾ\R�(~_?Y������K�q2�w�Y��;B����Ctc�c)�Z������O[(aX�ĝ��͘dC��jI��q�o~����ӲP>S�7}�Xm,98R�G��AdRP���Y���Pm�W�|������6��_W�Z�^`(C��B�*IxOuu�i5*Rb �k��[xrܕ"/�h��lj�r͏�T�\�YA"���[zw��g�Oݚ�>t��p�n��q~�d8X���,�#d��H��f��S(��`|�K��_����7�o����2BIh��$
ϲ0L�v�D]��"�B�i�z�˰Z��e(�O��`D%��f�_�{�uE�,��;	| Y �J�N������Fm1>�o�~�-�M��q:�{r�BÉ�g`�N��%�d��s�����!i֤�L1�q�}H�e��j��`C�I� 3}^��jO�i�xH*�Bk�];Sb�@�!���N�Jlغ��N���TA3�����Gɑ����Z��=M�&k`����Fj��P]4��B ����Yj�߃�vzh��H�t�5n�-��=N�\e�V4��q��̗:��D�������������ڟ�M���_����,r���xD�ɹ�l�}^y1M�XVv�U{�u�Hoos���ۄ��M����������� ]��bP��L��^�N�ydsn.���0h���꡷e����Io��~\�!l��{"�&�_"���lM����9+�8Ed�ꀲP1x�������G����wY|ꬢkNT�z�?
�l%����4��9Hm��:�(9XZ�ܖ[>�b�8��-��Ii�Л�K!�� ���a����#w�7^�q˕���k� b�i���<���ݑF��y�"�g�w����� Y�r�z ���=<9��%�z'���mRP���c¬�P�xgO�Qn6(_�Cu{mNd���g8Di�����onp�C���7� '�*��?��o�Z�5�cļ��b��;�Q�H��-�O1F��w��u��d3p���Bb�0!��	�������[8�褐�K���֤�+�0نcĐn�U��U�Ƃ$��R;�<X&q�� �I�Z/R��߶�Gr��f~���������j�ŖWF@so��B&���R�+���x'd�E����~�������|��%�LV�b�B8��l�~c!�B62���C�X�7���;�����-�/�a-�7���6Yܠ$��L�p}q|�+�kRx鄸�.xs�����n��H$��]!>��`������ؚ��f�,�D�|N%���cW��8��G�'���T�m8�&	N%K {Q>]�k�橌,&o��rC���RY!x��ie�Se��[~���|���:Q��m�����b��y�`)ه�r�{���NR��"2�� ���/�+�b�>H��R�6^N?VT�����|��ݲ=s�<��oP�(�V�0��:*N{�0��y�휃V<�r��2��M6S��g̝�\�_�]/5�S��׎+0�H�&}J;�;r]���C���=����r��W���m̷^UA�%��m��cr~#��1���;8� �TFQi)�'�V_�)��y?�,N^�&m�����mV�o�
EN�J�[��=|�e�FZD
������7��tr�Ƕ�Ge���բe�g�zL�C��"�B��<J.n��s/��g�ﱩ�J桵սP�De�����N��eZ���Z�cE����}���y��v�k*���������:�C��俖[ ��zc��ؗ*��3Ҟ��m�h�D�O]1�~}A�<���ߵ��/�q�OD�=^�a��&M���a6�\p/[�#|-Զ��JF���pJ�m�'g4J�ۖ�!��j�_���bTo����@ ���Ϡ��H�����;vo�7V��,���1��}�7E�h޹}7���e���{+N}����hhsH���27�A!1����H��n�D��"�N�i��H�9���f��?��F#����>�'i�|�.l���\��հԇ^׻IOB�ۧ����
�����<��uن�t�Vab��qP'��f+�3f��-d�.��@��xJ��!��!������@�훂�=r*���.�u� �8O�J��Hh��Ѿj�퉠vH�ef�_y�,��x5��9��UC�b;�^�M��`*z]`|��:�?w�$'�fm&�hH\Tu��&Cc��[�|X"�7�{��-*B4>q��)��]i3Q<�Pp��ں%���0���E|m��1
�,)t:v�m'p��v�J�ĳPdQ�R��f}�0���A~�p���?�H���+]���8s��ո�_%�tR2��Ez��C��$e� zѕ�V� �~:��r�"�'�u7����2�$����ʜ�)ߥiS�"
W��R-pt�t4#*}~�v��-�v���(1�����"O_;�<Qe��u����p���G�F-�϶ ��$�(���BrA�e�_��_���Z��=��E��)Y?z���|��:u��؂��[lhp=�.��6�~����_�"�w�ոX�H�İ��#����Z��^�_������G~���SG
�˕���� : ͽpmc������q>Q���e*�c�Y�ήb��&ﮪ�=�$��G@Qi\�l��is�Y$��NP/���(�q
%�#hc�%<��Z�ʮpf���{z�������������ۧ���lќj�+��.�mv��rU�H���'�Ԁ�[�抲�~�T�[?��'lǓ����"�o���69�(�#������SAt���ہX'���_[x_,�-��₮�g���X�叵���f��s�����:2�a:�����=�2��ա�ԛ0�c���B�vśR�Y�QA6L[	_,2'��S&� �T�+
mȣ$�����2��=y-$uRW��L9>���JW\�^ɩ黲��g�ŝ.�g�j�6ѭ�ۊz�"�Ep�-�h-���GS�ؓ��a����&�<��%�}�Zxm$ի>�4��<]"��V�T����>�ǰDX��P}�O���2�����v0F�(����@K/,�)�Y����*!(����YMu��!Kѳ��;f���t8�R�	�09P��Kqo%p4抾i�{tv��%BL�]Z}��i�\��q���ds,;zZ�ќZU�E�����˒���T�BO�$��e�.k��47z&��}�����Ǹ��dx�,�5�Ɓ��W��D�\�D���W8y�g*�~�=e|T�+P����@������odW82�r!:S�Ά6Hq��|mw(����;���&8��3�)�?���"Blr�К��$�/����y���y��hd�Ӎۨ�I�h�s쩗L������1��\(L�-R��oټ�f�n#�ɶ"Q�S�>l��Sm��O��ê�|���6�vi�!��bl��@���Ӯ�>����~ʶp���?�����Ά'���t�ːnG%2qӨ���I&*�^���J��y��(7���ϔ%��gQs�do�	����!r�:Uy�;��Iy4���z.zU����Ȧd�NͿ���~�T�u��"�8Ѵ��,��;҆��p����߈ȍ��u�S�}-�GPS��5�g�f�yg�f9�h�Y/�M,7�#���}1�QE��7�Z�5��T�Y���I�M�m�[k\�$g�T^�,q5wwTf?/��+�j\�E��h�� ~)~�hZ𢭝��11fGl�I����h��N�S/T=<$Ϗ���W�13�����3�����w�Ƶso� ������n!�2�C�a%�W� ZW��"Y��E�VB�����P���{ ع;ǯ��m�7G������)4Hɠ��'�yl��he���������hC(
;��?:��r��y�u��"ȓw1�%J�;�D���H��{T�Ҵ�\�1��OOf��=�Nz�[AٟS��~��?a�s��@�v�r|Oio3d���+�����H�˃��QjfE�E�U&��!rS��|�T��#�ɡG�jU�ªl 	�#*�E.S���4�~l�^rQi�׊S�p��zޑَ�?�e�｡��x�E��h���{�VDsB��M��8���v��[�l�1)�z:G�H|I��a<�h�
�r6��=��B�wh�t�)�\�F��������@5w{�Tm�M��LU�q�l�Im�%�"�Y��6aE���+��R�N��w����O��a�J�|(�2��o �X� 0A~�f4'b!�S�2�-�%C'Q9	&�I�(B��ҝ����k�7� �ڷ��bG�������{�uY���K����$��RV�����ΰ+���Q"��l�O~�w��T3�!�����%/��a�A����C���W�F��|���eWi]ezĂ�Gs]��ūm�r�~�ʰ煞���U����׋�BE u�����&*����p(e�{�II0R����7�^�i��<�[�( �{8�|����H��<�*�+�͌����K��;�P�H�z][&Hs�v�X-�t�^ey�Zf�k�`�K�f�MP�L�|��ؙO���h(��r\�o�(����oe:���u�&���~�C���^Oj��t��ROmڣ�����|���v�|n�OG����!LJ��aS��� �c"�cX֓窭!H���(���C"0�pz��ky��L�����^gSt�ݕh*��"� �O��j�E���,T���"T_8gH�P�p��-@��۽���fȉk+���c�:f�'��O���>h_�fk ��qW�ԩ
�i%"��3��F���!���Ú��gb��
�x"�'�J-є����3�;�;W
���m{�ΰJ��|�hi���'O��Xk
?�<NB���k�C�ljhe���M���ǝ�|�|�KlDm���u��J�Ԗȴ�� ����	��n�1�JI����Àƞ�C=�Ò�Z��}:հɨ�A=�+tJ��G��
 pH��E�5��"u�o�CP=j����x���ŝ+�1:��n����N����C��ϕA���b�~��VX\��K���WA��MPS�Si6U���z��C�o/lv)@zih/ɠ�C�?t̽�+Ա���<��P�j����}b�v/�۷=lkX�w�J�t-�"j�`��fq�p�ŰbuI��5&[�"�{�%�;�O�E_\0uU�e�<�����w>ۚ�F���S@�Xaa��%
�����%f��X���8m3T_�u�B��D��VJE� DUCz�!��CI5\�T��n��=vȾV
M�?���о�Dܦ]���%�=i���̣��!|�~%�z���@>�����;2���	�Z���;�L�\�3�c�O6��D�Ž�\�0�t:�s1��8�̦Kj�sB����'��4�#�Sx�u �6o �DԱN�J- ��H�J����J>#fyF�_?��6\�#�1A�U���ܟоD�}q�`h�ecdUs7J�L������(Ok.�1�-u�|�:��aJ�r,����y�����.�)-NVW�s!E����,��q�}�Qm��y�1��˻��}Q#���l>�/E;�&;I��LW��ǔ�ulMQ;�&�J�י��^�7L_�m�(O9��:�����%}G{���7i>H4;a�0��=̑.���v}������eBt"D4�$����O�� i��A,�Z���2�{�#6� �� U?��۰�܎>��`�  Q�3J?��ɒU�SKHr�$]���>`v�B��-�+�������STy�yO.������օ���4"���?��
������}�CpR�2��]$:�.�l�\�o7��g1_�g�Vbp�����R�j�つm��͢����b6̉����$���,������c�ʋX�,����`�qu5,�K7�e�~�G[�Z3Lխa�����.S��<�\��8�;�Xw�;sCAX� *.^p-dцq�N�`�;qL�bnʣ�����X֔�b?�ݕ��]�f$ee���+��" �۸��ȶ�.;�7(�p��uqZ����� x��;�W�,�(,@��BT���4���Fq1^��i��ʘ�Б�d�ō��~(o�|��]i���2��n����ˡQZ�R�=ʚ
�%{�>�������F�禝��
{��Z`�Z������hXG�0�\΂�~�F̖���
<5��
ʋ%��'w�L}%9���6uC�"6P��ǴN� -�ϙ�0�1����{����G��<;E};0HiC�/hs�aM���H��B`�P%"��:�D�[�w���3��,����Z7��R��Tn��27͇�Q!�.��?l"�
=�����;�3o�Υe0�0���fO�oE��3�����zb�gn�[��K�W��t�����}���ދ؜�j�n�nȅ4Ku�z�|�+�ӤӖ��e����T�O,��r�^�2�����I{�,���m��LA��.���]��	a.P�#!/T�>�|��Ubb0�����k��XD��^dw>Rj!sC$� �Д�e��������!�U���
R\���l��Ң"�nuz��)�t���%��s)p��?�\Я��g�Z�}y��
v��T^��%���ą�:�����I�$&��3�R��h68>	�_�?�}fH1{��r�Ah�*�Mc��8fM ��Z�C�8����-�*� ;�jpB�p7�*@ҥp��q4-ؔ1��/�U׉�κw�?ig�Mfm@���O��w�c㿶�3dF�������&��^�
6eUp��qd�=!�1􌒫�z�q� �B�@T��Y����Y�]4;�x����V��2"MC¥���d_��P�#��TD�����A�\F������F�Fig���Ě
¹�@�W�+��KD���|�w�J.tC�6h؁�%�*1��&�O,Ja�d�=��w�����|<�����Gy�o,��9�}�i�rh�����[yrQ:���S[���H1}t:Go�@����4�v���]�����1}k��	l�>w���9���3���6Ѭ��Q�]�K��T5��&DsǛ��e�Oc��� [�
q�^zl)���| (���Ȓ��_(�iZ��F��N�{�8?�Rn;]ع�~A[��k�d� ǪY��5k����מU6a��;~b�-�\���[�ƞ�'~H����8R��|%��2���PHR��Ta�
�7�XE���yH��h�P\&�����w����nn�k�X�"�����\��v��j��
p�0�8E��[�-�;���g_�m�g��{!��<r�)����f&#|��\|Q��I��H
� ��?�ob�O��1��I�mK�챳&�|%�z]�tR������i7U4r$�5�ϼX�Z���1�21S=$���B�� �05���A��Gm&�z#\���i�~ͣ���G���Q�&�D���_��=�%�.�|���~H�V(r���ר�����N:�y�6�b�2��?�㊜��>� ��?��G@G�¿;���:����2�|��0(��SS����g�bJ�2�M�XkC-CXzV
5�1�șO���e'�q$/[*_�pґ|-~{ۗ��jp~�Lrc�݂C��^��1��n	y�}��Vll��w�G[����,Q9㝉Nm���FH+�Irt�u����?N�5?�/le,�l�^�oU���4���S��)�\�H�ka�BAE=��:):�nv^@�5E����ǥ1��{-�xj|�"J��[y^�i�μ�Qq�\ފo6�%\�5
���n����O�9ͧ]?>A���r`�ltp��Ұ_�<:�<��k�^�]J?�����Z�Ul�*�u~v�uܫ�Ǖ4_�AS!��E+��B�����*�l���J�	Mj�|� ��� �ej�f�K�M_��~����8�ȮB�}��!�z�g"�Q�v�M++�z^&o���,��.�?���u�"!�=Ni�4��<2>��[����t����r'�E�5*f�쀅K��O�{gq�cgK�B�^%4X��&��5 �����~�h�Y ���55�))2qi�F�
k�(�G�L�NLM���2Dye��`r^��6�Ei��N���u��:���y5��8Ệ|��?e�����~�������ŬNZ�0��$���&i
F���k=Y�ye���4"I埱��Kr/���A���<4�+������%�|���<����K�����R/h@�f�O�6i��9&wn��Ba�S0K�4�{�g�������*�����/"i3�����WKÉx��+�D\2���d+��js9�|ƌ%��A}E�3~`�V��Ӝ��p^��N�[V�1&���4%#(��A`���@!�*=���a	{@!�YOi�(z��3�BԆ�N7��y��y�(�3��*���"F(�N�v�d6�*s *�C1�~-/�:���Gs�@5�%T��YC�f����*�BոN�x�I �q+6T��k6���f�Rd� ��T+�t��s�K���RM١�D�^��Ѹ-�Wt&*Ǎ����pN3_J4��ֹ�QO��DyH X��qj�q]�����[4�|H�`b�������H>zNdQ(��	^�3)P����d��WP��$Y��#vmO�ߖw�@�(z������s���	����Iޣ��^�)���Ԍٍbܼ.-��W�S�gN0-��U��K�X���D"6��՞����grEx)�8E̞�Z���U�NK0;-��vW$1̘Q9F /Tt`�T[I�mV12�d(T ۀ.r�j\�Fd�d(����f�C��7y�(�B~wT`Ho�,X*�5��1é�2RG6�Q(w�z	�v���N�:�׺�s�I�\�l�[�_��e)����-C�׍$;oS�}�T5���8W	��B�\UGgh�|؄������C3�#
̭�PoQ˜y�#�J~$��uy���j4�|Ϟ�o�h} ����'���:���߀c�L�H��#��Y�蚰��D~�KD���)�pД��0r�F���L���*�JJ��7�z�tH��޵�EFt��t]���D�=rr����c>	���n��+���Ή���;;w�^1���_�<|��K5K� GK��=��L_4xd{�(o(������߸+�&k�
�a�`����6�NR=}�qw-8�bC#��}gFa��'�^�(*��� �C�|����B�Em'�&�W���������b-��g�Ж7P�����ڭ�-�Pֻ�V�|{U�t �@�?g'{|\�3C�ǧ�s���~�0�4�b^$f��8��K���P�X0z��ق�����o߽�~����%*01�3�H�"9+S��dɥ.:�0)����.�1�<7|�1�J�g�Z�	�U@����~�*�q x�|`:��z<iB��b^�H��d�u8���VgM�)j��m��NdD)�+�����D�7@�7u���%'�~92��wϚ-�\��N��k��o
�`v������AT<M�+v��U���C��6�]�p��ϳ�8Y%��XI��+3|G�)��$�Ǚ�J�X�7!`���d�/���ռ(`®�5�.���-����G���y��7T����I~���e��hUG��nZ�N����jIR��x� ���c�����c�~9t�zR. a��q�}�(*�����V�٧�d��'�RIW���+5]Rd�n�R&V�~�����h=�w��X�ñ��,ߑqAnr^��<��}��fG�Ͼ���s4���o���k[��� 2����ZD"��v�A�0;J�Ъ�d3>�Z��V�	%�l�W�pt1j���
��Aȯ�i;2�c�f�ʠ/Q��XxL>���,~�`Q��� :ѨR�����N:Y�[A C�=�$��w*{�?{B�	F�&)�
\+�j3�Ȗ��kY��m�H��<�ӥ7���G�_G
��9x�"��@4�-g��2P�GFG����5�]=݅B�?��
l���{�!Q��g��
�ϜւC�r�Al7��OB���SB��q��]V'�Hz���J�$i%M�!h�4��֢���z �)Q0���YJ�D(Vɾo>�
���L:ȎA�h+��9�E�	��UؚX���bXٳR�[��	U\����L����4J1��4�baHl�,��nS�����PU���hM�N��,����Sc�rP�b��(i�U zq;()���Y�[�'̀�Q3m�����Ԩ'8�TQ[�����@�K퓮Q�bC%�5�+!]YU� L�;�ͥM�f ��(dZ1;��a��4���Y=���AS�1�%���y��S�����@}pC��+G+��vq�tE��\AOAC�:T�??eK}��N_܂����!��  �]l��k@*%ȸ�`\0P�U:ޖ����x��ܠ�8;-
X��"k;�?��M���`HJ�]���Q�T��S��G~������JR�8��
_gvWhg�������Чټ7�>__z�����v�d��}$r��er�]��&�փv|й�V-];����Wx�W|�ԴZ��B�A�a�u+%><��͵���+�7�S�!�w�Vt>Q}֒\�.yp�,������f��Tb��-N�����,Uevh�G�9~�3[�L�|_�N���j�op���jX�K��!����_� ���p�PQ��b�(;!CN�f��0Oչ����Wz��	���V\Loc�.�}��W�0��P������#��
��c�[6��	$�q�!� �~}��K�H�7x����f3:�`��,kV��%� ����o;
�]L��U�
#*p�q�J�Kz���qD�on]os��g(O�/+�=��|�7K�]�\�gQ+�l.p�]O��`ZE-!kM��Z 3�!��L!P%%�*CY�J�?�� ��7��D%�f�ҕl�Ppʹ�	u~�� _�*��S�B=��q	X]�e�]�M��ot���XT~������3�BF� [�F:܄@sl>S�M�K���Oa�&ia;��sM��w{8��/{f�影� ���@#<z�-k�W�1�wac�DtرD��KU��z��k�W�Yv3� Fъ����`VY^ϴ���>(�?7��8O�b�tӜC�ոtb+e�a�i*XfJ�U#�x�7E��@�ک�����x�F���p�4�7b��5P:�7�X���֣\^�#VM���ej}|W��Yg4'�Rڷ��#�)Ǻ�>1�C9d��)5����R�N�qTץE�64̲���FՐ3וat�D���=��-��#���H"�u
84�\��t 66P`p�ƹ��T�;�Z&��T������.�Do�銵/�5��(�]a��z�n��h;�.���b�`?_��% �rWGs�}�z��b[�����̏�>��ofWy9}b�3(�z�o���-�{��]J��,��/|�c�Ղ�������W�2�ۨ[9�X+�ӟ?�H��y��������ă���Y����DB��VE9R���5�Ф|�#i�A���ȕ�L�ޥ�� ��E��ZA�b7��m�K�ª8�^��,�@��b�"LT�%���=r!W���d���;��	!z(�e��2��M�P�xfw����𳨽q��f���l��!Yf�a�pƂb�}HJy�b#x��s��h�5	Z+�R�d3�/�c��u��	W�ph��*9'F��E���)�t�Cӗ�饺�Jz$�}���w�Ь�����{ N����hi �K�r�	Z �e�2�����}AHШ'��Bi�[�d�+�d���_D�V-E�ɓ6�t[<xs�������_Mul	#*�c�˄h�����Zb׬#i%�^\=�����[.��an��8��C��O���ц�d&�Ť�(w����#����`��]�ĺG���G7����b^��63�s�WM�SW�Y`�aoR"��_n$Oĸ�� �Ŷk��|d�f�6(��D�Sw@j��r�)>
Ǫ���;���T�$i)��$)d����{�,��������%�����RM���}�g�OH�7�k�\-X�y���n���0Y�������EN�۲���nڋa�q��H�b����:�!ؕ�?�%8�b ��4���[�JG�����}����9N�/3��&�.V�2͂�B�YQ���I�mE�I�g���}@�*A���4m��IY��w��R�:���,z`�T�k�G���zeG�},�G1q��Փ_��ґYi�	��3E�0 Q�k}z��Y�E���9JX����H(�g7�iy3��(�S�1`߬[Ͻ֐á��^�.�5�[��Dy�C��^F]E=��ԫk ���ܠ���31s�S�����zB��
��8,a0l����C��$w�o�a�R:=�xТna�x���3_��@�;֬��T�s��%_ Q�S�r�bm�9����I�IGٍ����r!��;/�yp
[R5�,]O��O_���|��&WhY#�#�HS_3u��烙���s���V�{A� -2��ڥB��S-�C��Z��Ѳ��pO�>�3�M���#�Rj-�E�*�<!��
t��V��#�s;���V��P/�7�%<��s#�3���PWP���P�6ELv�F��-����@E6v
j�dҖ��­ddz+@�V�z�*�~�0�T�"���Q:�)Hx�l��=�+�/Zg����<r�W�^�~�����w15|q*`���(f�Ž�;<�%�m�LU��-��]�O�
���kڲ�=�,��24��:����>�1J@��6\J�Lޕš~�����0@��3��Tyr�Ш�� ߍ�p΋��/�i����uu�f���C%�?5c�YS�.����q��O�^ƢU�G�#9��q	��
�l7ĺ�*V{\l���*�l{���qj'�Ȣ��~���O_ɕE�o�g�>�	����EB�|=��$�G���u"��:��\4V�L�tl/5��O��q֒aǠ���B���5tJ��9���V�{��hQ�/Ǖc0���B#	�!����Z�k����������yq���b�;2C���6����7_[��������7�g�Q�s��h�Eh��L�iwEN��3��}O�W��2���C�ߵR��¨ 8!����Ү
�f����p ��up�b�4a��4��0!��aZ��;	�X�=��b�7e#������b��lt M~C�b �9%}}+������
�$�E29���E��1����L@�[�=Gj|�
�D$^ �μ1��:�j��ƋZ�$�Mr�2�t�ɫ���-p,���u5r������Ƙ��I]�Q"%����s��u�r�������F?�y<�aQ����L{��+ˁ!����g��m�A�?���>ɥ��5o����Ev�rSi���j�/�Z
��哔'��7�~�P�3��4�c�Q8U��[ѱ�>�]���R ��1��? �Q���֌��I��E�p�N'���-`�P繓�o#��_̥H~vt��7eLPN��&��s�Q�_�m�䮺S�=M^�梞�Z����W�ʳ�-8�J�Jk�q/�q 1?x��,�A���|�_�V���Q�x..�7�(��/���#v;�B���]���X�/~R����%%�o�����'iP����7��H�z�k1��hO[L���0,
��Y���p�*� �)u�����h_)��H�R���@���P�#���2$���YOI�m�^�����"9�@y�,�/���E ��r�*2m�/�X�/ljý�*u���	ޯ��D����A/R�I����6��`~�����y�%�b�}����}q�JC��Դ��z(�w���"��Ly'�4�$���.=;1S��l��\38�cS���̈�FxV^کI�,�9'��I(C<J�L��m��[��uu����� Vxv���� p��UFgCv`,���e^+��.o���@�뷳y�?���x���2����e%�^�dt�@�H�",�t���9cM�*���|����+yk���ڍ���T�"r;(��W�~\ܣ�@b��C۠�h�����#���6�.w~_%�eAQ#l�M��}�UY���Ϲ�
;r�B���!0{��5��` ��-���Ku�r�{ v��/ w���7n�w��7�$X�n0+T�h���OZ��9���}��?�L��w�^��M���,,M�X�¼Ad)��v}�Q�{��&3�q5����XWl�����~���Mg����$j�m�:�'4�hRy��^��>��#�y͢�)�����-�2H�D�8�m*sn��A�0��P�̘��kE���,i������x��F�����j0�n�H�\����nc�(v�����n�}��t���5Ֆp�X<w���Mm�=�n��Q���0�HՍw2��q]�m9+QH�fݾ>@�*����qfS9^��R;��8U���m�j��^�@��^Tɾ���f���|�?��.m����X�����h��k�7���2V��\��y�-����ƅ79���3c
���Yu����w�#7�YC�,�h��+�E%
 �܁wD�Da���{1�
�}�<6+ -g�p �S��B�|(�qKS�������My�h��Le���Yʾi�/���ag���@Xkި��A7�����`ot�EO�H�0�-��3
҆��$��5ݏb%c�DK��T�&�ڔnhl.�Q��.�sp1,y첝;�JKz�>ɛ@	�@s����2+�Cq5�Qz�"G
���G;��.���bu0*���;�(����� ���^��줍�{��e���㬃��s~��'��V䛇D�]�R<v/q�+-Y^A?�DK�Q#G�m�Jf�qyôW��HVR�!���+{��E�(N�ѕqсz�9�+	���o����U��{���_���w\���=J������i�+�e*����J:@�.�,/I�9�y��>��bK5�A�'��t6$eu8e�j�o����]p�I{ۛݻ�}9Y�K�.����G}��X��Ҏ��d�MKI�/Kc=�(��.�}k���ז[�o�:���G��V&2��� ����A���ec	qVsC���5��h��`J�-̊/$�,��"mKi�D���d�I�d`�jK+�n�g<W����_�+-�߭�	���>q��ּ�c�
��To�<�3xEiK��[��%T@I�Io���͗]����m�_݉jy$����C?�.�Բ�/F�x�6t�Z�fG���n�A�WE�<�$W�v��>*�	.��6�H�R7�>��&ݳp��;��+�:YY1 5��x���� &�}za�^s̀1�`�y$��C���۳<��/�a�U�X���K*����*"��6�1�3r���w��E?�R3~*I4�G�%X���2���͠��30l�k��ä ��ꄌ�}C�/M���ZQM|�{��Y�7�b�K4��(��t� �,��+��!��靶��
�a��λ4���{�̀*Zh�t�����#	t3H��'4�����e����L��Z��/�z�j�a��|�>�����Vʥ5���+e���zS��V�=�^ߺ���!~Z������A�.�"�\@��j!�j��:����Am�a�8m���9���x1���:>%�1�)�~Z)�C"��v�S���V��� @��Yc{+5���룸m��^��h"%0��uo�y�j4�p�g8�sV![����+=$8?�'�]�b� bkk7��hV.N��^�lġ�d��7��YO*z���4�w@T:�#L:��fna�F��O���?�g�����'��|�;sV!W�J@~�3�m�����r�0���B��#x�ͨ0�Eg�����6��e0Y��%y?�R�)�P��Q5w���NH�3s1o����(d����}�_2H�6�����,��p�ZCH�J���ݤ��ӱ y�Bڞ!(��]Ȇ��7&κ��O�w@�uA�S�3��w����1:���W�q#�輴� �v����9إ�d�]�n�s�ѿ��=�>� č��y�Z%"4۫e˫�˕�`%7�a�2����d�Zy���ƾ�HM�K�jV��kw;�,^_��,Cd&#.l�-y	m����$��)�a����Q=��@h(�m�P��8
��MuT�}�#��8QR���}-�W-?�Qg�:�m�XC�k �r0�� �hd�1��4�ؼ���`�͍�N���Ƹx�,�>Eq�Վ���3���·�c{7�I�~��ъXH�"D!w"�������8ݘ�R��m��[�jxd�)��&��'q�ߊ�.S�!��]@���;P[�A��j3F㹧��8Wb*bC�1�6t�;�9H� j��� ������  �s�LP�6:�j[GW��O"�$��W�PK��Y'�b@B�=�2c��O�	V�'�馶�G���Uu�������~���� �ȃ�)n�g�q��K{2����0S�4���eeU�ߍ(��e�7.�����&^ZZH��V🕌������+oO���uŗ�n��J��}��j�ߵ�wė����(y�h5��"���eg��X��/��@�^-ѿ���BV  �q�t%{$�0\���8�564Ǥh�bq�#N5��<���(� ������3L�υ�ȠV$�D���S��-ז�{9�ݨY5��a�1��fA��W�T������8Bg�:>�.�m�""EbQ�R��t��W���8�=�1���&����X�zu�����y���	��Aw"�-)��6�Qv�"U[é���j����/?؍�m��Ȕ��F���n�2(Q9���9j��jg �;��Ď�tHwSbI����6��?�EP���a,A�Pu������ڋ�(��3t,��tk� 3L�@@�['��Eg��3�"��p
�����٫��R�n~p��o�w�c�A]"�č8���||���K5!�2��wNõ�����u\s΋Llݾx�QM"�% &�h���������y<���ݱP�=���46�<�$s�C�R�y��݇��O/��L�w�I�NpqU�W����3��ZCR"
�@e�Q(z�y�O�*�r���آ��ZV��#�Q��K�G��2�q- U��;�nlB���s���G�3q3�1W�^��?U9&�K��.	�m��ph���si�?w���%�S-������v��/���2��G��g�t����V0���x�{��*
��~�NX�VtpZ���Yf�9̴DM�GE�$�*蘻�|�z��1��<'�!М7-.��u�=L��;���nx���CS���T3�Hp���#J�j�n�
�=3�D�:1���	Q��*RO�0��k�(�R��m���M�,r�:�$�0�����|g�V#��\���?���]�zeK��V)�5pA�6W�&���w�IS��2�'�"����L����P��"7bHLa�����v�6L�:50N:��im�S6�0�64 ?�I�8ۿ��`񊢐��#�J� ��b~r�n�h)tv�ٛ�����=�v�C������,�6�n�4;�W���lvo-ѫs�w���>�l�<���&9= �M�5o����F�������#���}���Xq���-��V���!�Ί�$Xh�#�ώ�p��a�Q� s�%�FpM�:q�6��WI����^lj������\�2���Bh�z�GL�ky
,~εB�]���{��ks���X٦�R��&J�đQ�xعf�e���"�`4�.�F���ۅ����s�t��L»�J�&�����w��D��_M�r�Lw��U�S�;����R�yv
�<LX�?��\�7���{m�OW�d��>E��w��K$�p~JR,��d�����&�L"�h�OO��-�)���<V[���l	91-I3�w9����Aꔏ�ڔ��nw�Z��P1N������ Q1$�'9^0y�2�)YL�3�?��*���3R��TQd��8����%Y�	��a�$����'8߾0����C��f8>:9�L�P���&�Cf|-���h3�V��=���o�?����r�z.�ua ����T�F��� D�4Eo�C���h����k,�N�7S8��v�׀]�w�r���-�-6�zꙔo��h�fcbJ� ����J������#���$���%��F��h:���Wdb]�n�v�-ӂP_?��7rQ:�v�S8LWJ�����Iv�
�}�%�[ќ�	��OaHA���R���r���R'ap!@A��k������|��r�A%�at$��q:�E��Q���'y�AG����� ~Y6�ۧ�!g�Bg)����K�@.Fw�%�L�tĻ��R�T`��a"ڋ�<���R���5�`n��*<���hF����^��C���z�rxc:PBۛ+�3Q����B��=��rU[;�"<��K}N�y���#mび��Vb�����n,P��I������>���h���M�/�������T�Δ'��g������kqJ����Gf߮��\I�	B�񲀿�SP���$�ED~�V�0�f�IY��X�S�RZ��~l%�4��7!���w��)o]�����Q�?#�
�ug��b��������D�#mM�\ )�F�nF�S$�X���k kv����'�{ �~��]�w{)���,��l�|$R��-�8�ُ��j <��"�S��і�Hl_�1!�#)�)��x��U�:ߞ@���)df@�Pm��8fQj��t�/I��mP{%_ǟ�j�|Tu#X̡٭�p��J�L�@ۍWg�I��\y?��jW�ܡ�v���5@�Hq<R�Y��NX�d���TA�迣b[ٵk�(�(�%���Ȼɫ��T慛O����ꖦ�?ۋ�2H�<Y�W�?&��Q�*%�v֠y7!�S�![�0���HX^��@�����	���z>'�/>s۱�$7L�/Yv����08���܋�eX�L�<^�?�Q|_�1Г����8�%ȳ_ܦJ��j��Cdq�˂��M�5峡��HYv�Y��(�&�ध��c���^�non��@KK]\Xj����UP���t��}������W�w�(iT\S
��qc�RsR��X��'x312%�۵��c$N���Kxۅ��Q˧L6e��2�Ų0�����-���J��"o�'�#ͭ��G��SWa�\1-��;$����������*Cւv�(���;����ۣ��/��S������8����9x�M0rD-g<WC�`	[��(��͋Eu8>�sv�T�{Hፄ��n+�����zO_Y)�Z
o�>�4���Ma��k��y��c+IB	�`����A���"y�w�DR��	k[&��H�h�Q� �'n��۩��±�K�9�����7�!`Մ>���/8_�n:���g4�+Ô���d(I:�z8M���3dM���G+�o��$�wʌ�5��G5i��H%4C��"����ߍ�F(�m4�d�0�n��J�Y��Ø�'��Y.1
M�LCt�݋�}���|��L�S{-%����mx9������Kڦڒ6%���o�?C����������N}�^��wq�| ����3ܐO��m�3�ы*a0Հ풅�;���z�ם|���l���Y��s�'P뚢���E(��wQO�i�/
�L�H(\~x� ���>r0L>;T1�W4�X��M�^
�wc_q����� �X�^��v�AG��-�9\�_��yէ�����e�pr5D��h��껎R��}s��.I�<_�Ŗ(��پ$�­Kz��~�?CK4�oC��/�֓�-�tE�Y��2�et��T���%6͂H�'(��\@�)�:8��Ni,��p=!����ٗFiF�(�^�;:yT�/��QMO|j��n\������|%@�VЇB.���c~.����@*쁛��ś��>ߺs��Q�*�K9ҭ�u���c1 c�A:�}+7P-t�[X[��F�Q����]�}�4�����s�d'�,K4(� ��ξ⸠���mV�ܶ���&/u N(U��B��.��a?�c�|F��1��=�\��fʌD�|���h����YdI)ټܜu�[���w� �y������G�J�u�w97娃�n9���6d���뾤D��[y&D����둲D�j�Xj�:yq��۹��tJ�-�:���Nw6���mZ�.;2��BR;�p��@s����n��DU��5��R�����.��F� g��2��4��7b?�s� ^*�P�[�0t
�ϾN�qE�j.�{��v�U�I<�T[� k��_g�d!���x=D%�GeMypu����ӯ��4,l��PL�o_<�iP=�UM��,��o�@�B�_Dgpۚ�j��1���,ŀ�t[HE�ʨ�����$,�Q��!��T�1�����P'���r��b2:��E�ɚ'��'H�#������|o�Z�����Zфq�ƶ�2��͜���aڸ�ވ�r�,�Gc�ڎ�f�a*�q��V|/8��I�����r'�����B��|Ψ��O9��5�����;ˏ�b�Pw'��T視��� \�]���Yq"6��$��� +��44�V�b3����M�ٯ���
R	���_�R��0�:޴�*(�Tt�D�J	Z��W'�J���-�Cy����mԨ��^���GL�G�곁�܉�~	&�Y���\�E�S�0Nk`0�B�v�ڱ��jdP�oвh�-5����	o;�6��Vx?qbsv��ݔ��:+	�vT^������o�_ưtP�Z��DR�Aj���� .:R}+4o���z���&�&�L�F
y��>�o�V7&Z�* ��q��C-z���~��	}P�ak�.U���
ր�|�#Q�V�7�eW���
쓷��bACF�%��3�QKw�:|Ѥ���K�@:>׫������1��q�	��SJ�s&�,*~�ә-���(��?�q�0����k"�Y �۰���2?�P���/^ԉ�i�x����ƿ���])
���l��{à��ݓ�Ii[Ll �>�M���\�bF��j�#�x�0��F�,<%�\f�R���˺ ��9Y0��qjk]J�	.���m���6ͳc�B#���$E��qq��܂�(�rp4��O��>HNl��v$`������ske[�H&�r���
��٤t�6�;���NT/^r��!�!$�
X��^9��߅d�%ھo!��ےW�g�z�[O�R���[����!����=�έKe�ju.��� ���"�4Ż)+"�����6��Z�U�E���O�V��+�3�ex���=�6�(,�B޾��%ΰ-�������O�y<�+ }4�z��D[��t�)g�c^��r��*40�}��U �at��b�;_7`�(�v��.`��A�1E&�@���8 �~�e"[	�m͏lg&������z���m�zW!�#
���������D�2�&uQ���U}P��!T�n���E���8�@H��&�^�}��)�*�� �B�Ҝ��N��&�*��N9�Ϡ��w�m��Ks/�
��R¤Օa�� �%?�&R�����/֐��PZ�o5����K��2H��K!�j5w��"e�"��	ܞD)7r~ CH�������� �郦X���	DK�a���*uV3}*��g�T&�"�/�X�$�.^sg\=J��%6Lc[2�3p鹟�����u�1[Cl?V&(4vf�&o1r�-#[CǤ�&h�p��O���t����O�7k�G�	�-X���,�7_����"˧�>If��sR����?ʺ��HQ_�-��F2��H%u_�4�!� �	?Ύ���VMعTH����	*=��/�
ho���*r�a��؎
Y9���(��w��#����b���B�#�т�w+N��^	���w�Χ�
lh�}���;R#�����	��VIk� �+��z��m�����j1��R2¥���������+we����
���9���K�wZY���gq�(NA�S+_�ʤn(k؅���pD&r�t�!�H���� 'c���c����]����si�F#��<<�
w*�+nhN�"Zfg��!�_�q-�@��y1�"�[n26�@G�RE��$Hx�%A`��{�ƖPJ3��շ����F�����҂`�D��Z��q���C ��j�@��F�C5��;#}l��������im1|�:�Vd�OKN �A�����ۏ.P��J����4I�����t/:��0i�i.�����Q�2�����H�O�Ϝ*\%�l>����Rw������^l�=	��G�q��F�+[O�>"b����!�J��*u���z�B�6#b�� ���F���rO�!mi��TF�г'��4�
J�<\����"  Y+��:%Ap���~ܐ]� ���2���N1?�kNn�:5�L��-���E�2@_\ KC�����-Z��^��G}�}2������PY�6�o�,�����E�;ru�.o�㡊$�C1�w�I���I�T��u.M�g��7�u�����V�I�-�0�!=�[`��v����g �K, �&��,��WޚH��3����स�,(�}��j�ϖ!3O��*�<��`�(����!��6r���0�X��`sɠ���Hv���aP+�W�u>.x:�6�Px�ǊUEx0������;U4<�{�1��e��:C/!���MJ�0�Ot��
>�F�!zv������iT(�������Y����9��:���gz�L�����d	��#9����V��-�&��Zn�?�]��s�=�0(~m)��b�$?N)D�w���On;��j�}�����wg��3}��(H�k��=��V��!�Xђ�g曮�_�&���T�}�KA�m������w���e��د����/�f�j�+3&��%�
lF{ɚ�Ew�K=�lE����s8KP=�.v?�(S
k���r�ڝ���_�Ҿ�Q G��r�V�4�����U`�}	!��So��U`FI��	�f�VV��y�<@�BxN�Y�|ܞs��e��_��(�Y �*  |_�l���$�f�Ho�('���ʉ�5?5h�F�5��e�~C�z���ʳMHb�_aG��1?�?�N�+]ԫ�e�������Sa�/!��s�`	���T�~��$���9�������v�a�K�x�49���Lҵ?֕ڴ�H����>
L<�ڡ�-����mv� C�j
�@S���/��&����ߚȲi���כ�?�����Ls���Ext(z&�%h��bғnS��69���_{��#��$SP�W�8����/�TO�
�'A�HD?z�h3�,U�ac��hp-�`M�Z<>3��\�Z�'I�K�9�H	d҇ �rY
Gƚ����"
�z2�����P��x���J�[	gr�����r}�Y��N ���U8r�����F���3�=�����Eޟ��DI��b�n�����2��4x��ѵ�GH�A��啪$��٦�0[M�UU�e҉8��I+����pl�O���t��W�R�a��_z��e�ǻ�� 2��1@쇇���2R�mw*�CнK�@l�Z�-�OV(�7���rč�����������hlg�.�C�g���Δ�b+�'�H�~��'d�<�팺6W��ªN)JA�v�$��^~����_|�N�����Fl1�?Y�ĩ0��q[�YƁ��G��d��0,�{{$e$���2�^�*���"6q��ZK*N;��� ��;6��;n/��hI�P�j�P�|@�U�r6c�.���ad��c��k��{��`���%D�T��kY���[|��&4k��c��;e��%
ƚ^&L;Y����\��+�ix�A����:Z��5��|�2TΜPX��癹ӓ�	l0a��篝� �[P�uSAI���2	Īd����fH!:)�
&zU��/c��$�������I1g�9R>��綨;0c/�1��������X<k'0��_BU��ō�Gy�b�;�Y��Q�l5�"��p�2��L���zF`���qf(V̈́ß���*?+�eHJ�j�R��7�ԝ���RR����8w���eWx�<��� �7����"�UGO�j�A������CLk� �m�s��Z��b�û@oS7�>-Òe�&S��� H�<@}4�}>ti1�/|�|�&K���?���ie������0FGW��O����噁(%��z�:CV�,H+� ��U�õ��2�~l��ޑOܜ|�f*��j;�ܐ��.bV�G�8+��J���o����{��FEb{��b׊��F��
(�T�U����'���گ,8,���|�.q�,��D��]Ip�r�r�}���MmJ��b�dx�=��D���}������5&C~/k�X����~�-��B���_+�x
����/�qk%���/�3=C�O�"�!uV�ؼ��TV��(4��O�S�������_�
�үG�k��U��(��=��W�s�ɕ��:��j�)��o2���r��ψ9����vp��})�`��q@���/�r5{_��ư	�ZFW��DSjA��5�OȠx�����>d؁&�`T�u�.��x�N^@�9����M;עgI�.(/�U�yU���/k��n�s�3b��)�<qb8��҆7��C�gF�Ʀ~�n�����aC�~�E�2D����^Q�ڶX	�bX�k���K8��?����駭g���%T���5.3)����������b��)CR�eo�PaK���~S|���hiz��?v��p�"��3�R?WX��%�����A���K���XR]���H�j���V�h�L�
-I�����<�l�4�W�:4��S��Q�H���7_`�n�w�O?�Sv��6im��8�ic�`S�m��T��3��1�'��~�R�F��z^��:@W�+����3�7��W~z�~���it�p	��z���m���?J���l��"��ܺ�gR�<���r�4Xf��F��9ֈJ�|�����V�7��/u���@eN��dz��ꈫ;��3��s
�v p\�5�?�nz�� �)�U�pW���Y%ko��(%.;^��"�1Nwʭn>.Ef[?��D��8��.��`1���V�>y����>���z�ږ7qF8��]H4#/��&;&�%
3k�RLg$�j�(��4:������/o�}�G�0��5R�����e�۱t([��̳kA��<�I� �=��E�`�CxQ��_��X�m��3�w��,�0�'���
���cڏd�Ұ�lA��v��f�p+�;I��^��a��,icV�?kF���`Αr=U�"Yp`�-�\u����/o��-�
����?�4<�~��x�ΰ��)�Q����2(� ^4�(&PFGݗ���_���U1�'�k�G�Ii]���N�g!�!H�}O���Өc[�q#��̦w���*������H��� Lp.Z�Oa<4ۆ����1?��q�*i�=�Ɓ����&���暇47I�\���Y?�L�Ͱ�;OJ�����������U���ŽC
�=^����9��(�;�熫}�+e/Cn�O���:�Y�n�f�r]�%��D��X�����?�^��]sGd��w�a:��M*�;�ٓ���>�U=��������FW�n/X�1�a�
�nY�"��Am�mc[<OH�
z�i�w��k�K�4K�Vu%A@d�9�5 g36k�_�Z	-��&G�k��	�`M�%�jh`�j�?��r0?���D��!r\a��R\��ǴǮ%��YX�G+=���~/o�e	��Q�̕a�~�s�F���>��A:�ʌ7�vnB�pߞR���%k��6g�_J�Tڠ�K�x]��	�*q`R"'����0*���'[#8�)�Y���ѣ#��t��p�V���v�U���z�{i=&���K�aO}ؒ(�;U;�/��/�2�21�����I���� *Q�k������{T�*������;�m������O�y�7�b[������&~H�D��>�^o�a���M��$q��{�3Gg<]q���{=����5&�?�wdQ��n�Q˒��%�#������=>��"��ΗLKF��pg�^�p��o�.���~�n����'�;���9Q�C�RV���X���4�],`UY�}�n0s/�<�I�,r����r��� �����l�3�O��w��W�/�(���<9��/8{������pRױ�2�.Ә�߿�dS_8��pV�
ztׄ�RIS��u�Kz�j�U#��A�䅋:���n}�(뾶l%mO��/^��8��h��$�&՝W�Jm2�k��Ujc1�s�g�����Df��a�����y݈$GQ��D�/@�ո�To�3<k5���'��$2L%��7\�g1��"��d�7��G^����0M��6�H�l^I�K�Ke�a!�lU�2N�3�w��Ccn�����%��FZ>��v�FL��#'+�`d��B�>�	��Os�|��2�.��ǫ53�fw":�/|�o'�m�b�]K/�Z}*�C���V���Q>�Y�` ?8�&g�1��<M��7R� ot��`��o�Wm��F��o)�r�I��?09  �Ɵ��@�{���nIִߙހ�*���;u�Iet�Q�<��������_�.�J�it��n��˨؆}��y��
�i�|Ǒ��ve_�o�W��=d�/�m@,Q���8���s���΅b0��i�(�ts��-vf�R�J>��$D�L���oy>Ӎ�FFtd�����w����?PEԑkX?r�'�&�]Ь�y��4�J�i�Y���'Q���'s�ZM�a�^w���I����吏����,�� ����@`�r�vP,��D�u��%�i�}4��[=F��|�Oe��xizmhDki�/cP�p����c��c!̌�E�JP�Wo���?���_j��+�&Q�؇��L��,^7d����N7�x�'qb��6��z�kp��_qy���YWB�BoH�<�rZk���I��Y�RcW>�(-w�]{���c���6_/�=��a9Ҵ�)�8e-K��yノ��֨J&����@�Cݴ������X�}GE`�6�d��7�\���N���c[���� �w��l�� ��9U��W���*IAH.<V[��I� y B�"�Y{dV;�	Kt�Ȏ�{yn�; ��[�DF��&�n�O���У��}���¸�1�����	Q*�sG��P�4������	�c�~y��EF��W݈�H�,���@-n�0X
tW�îBqY�[�XsV� ����F�tc�>HqI|q��"���,��3�ҽ]�����m�0F��,eT���aȧ���I��m�S�Jؓ_�^Q�%�6F��C'�gړ�TC�䐩Z��A~���dR�rv�&�X��X�������>��=٩��W9+hޙq�R���Ј���;[|�*%��-v4��j�hK��b�f2>nj��7 ��Na�\<\o��4a6^X����ȷ:GGY��V'㱇�]��=�����o� _<��0�^�0H��t?^c�i�`fx]���_����ʨ���U�0�2�p��jcY,V*�^���E�FIV�/�+���stV/Jj��G������ȓ���;�Q������l��ǫkx���b���~��.��Z�p��`.�q��>{��=�O�
�ɫD@ۘ2��D�:�J�0�y<*�z���$g�)�n~�cZN�l\A���ɕ�����MQ���|>�b���@r=
���_�v�8|oȝ�r���\O�!��+��B(A�$��������� ��q���{����1���k{�"��=�o?W�M����3�^��݁ky����X
8�J���zXN}PGL�C�{��o\���Z�F;U!taR��)4zW���+�{�Ǖ���q��z��!��РQ_���'C��;��SS��ҮQ��%[�c��}�P�#q�&������e�TG,nZ�`vʃ��Mh�5�]3��o�Z�k0~���.�7�2�?�^:��U��d�$A�������)�7d�go���N�͡�
#�;�i��ƴ7�w���]>��6s�r�X��ܰ)�%	P��7i�ɜr��!������?�܅�luh!0��Q'�h���JO}��`�(�idd5x"oX.�ԘY˽q�ؚU��du�A�s\`M&z����v ���ur裳��~�O�*~>��-F�5�����j�໬�sS��Ń�q:�L�ˇ�V���e��P�ׅ.D�H�{U�ϢU	!ZM���U�/5i�Y��)�3�������$��Xn����V^y�~��ɋ6GqC�6V�U�&(w~����\迦p�Y;,�eZꦌ�QM-&�Ц�ƹ��)Ip��տ�"Ha$��nݨ�N(�y�`��e��R�
��������Um�=[��kd�~~O��*YB1�=�b�"�o�gVY���� ��r�U�Fn'eWx�I������P�
0*O�j���7(Q%]�>�O��W:��x�PΠ���9���
P�[FO4c�Ʈ{)�E�򮌭݉���	1q���aq4φŦ���7W��s�`����ko�X��G�8w��X�H1�:��c�1W׷`���B�vtqdiЂX��qS������Ɲaz�0�	�P�z�ĸ��'�M���3r���	Yn
f73P��~��v�|�!p6��|�Z������B���-F��9��?*��r-�q �WBq��o��Xr*���Z�ץ*���o��\p{%�z�;��IgTi\��� �KЃ^���"f��fϝ�jAd�o,�,�K��4[�����Y`3S�L�<�fP���R�!�&օ��m[?;V_xg���֎��W����P0�����&�\��.��}�`�C�S�Q_һjy9'�X��Yt���CR(	�keT~ \O-g�-ʍ�8�T}��3�c��bp5��U��$><f}�A*�+YD�wO�����4��'��-`UU1��\�VMe}in�뱄���XM��-�W���BUw�{�zy�]���A���>5��f����ٹ�u��cHYW}�c26����v�/uş�jʵ����Y}e�D 3_���g�tw<˺�we�q>@�,g���nqm:��X��2T����=�n��O-{h�α�S� �饶u(�B��<����Zq�ĺ�k�c|XB����;ydl��^�
�ы��8S-]�|�΂r�� �Qe���bF6������������}vh�\8��I�d����^���/�26Y xᠹ������4l��L(�Q�v�?�	v�C$�M���9�Cx�����K4��A�`4��ؗ�x|���U���j����!'���T��m�������Btm<��O3�+�1lE�٥`v�S�-%�\8��pn�c�D),���u�%o{�U!�::P���G�P��a��kf�µV^�V�� k��]k�KP�0����ey��2�'(V:�
R98iU�@pK���R'�'Wh!3���
�[��Ff�[<��[��F�|j6��d�l���.,S�9^3��	�}��$�j��LD� �6�I�H���-�g̓&�(�Io�*��U�	��:��w�IA��81���k���z�j(��sjΛ�V���˔B���U�v\�M���`2m[C$0�['�O#>6���N۞#��+�ܬ�o�scm;:���19(�>ӣmpL��R����jz6�(4Si��n3^l���p���`�T7�o�d."=Ҕ�%窀xg�����o3v���9��X:�WeԪ+��Y�փ�\����_)�L�s6п
��kH�����-\]d�AC�����nh�B3��$���=J趐����}X���u�܌v���Q�eɽ��d��ǂ�0"�1).��x+��w�����������E>�b�5T1	̕k�1@�N��+,r�!ʔ���xpc�y�d]!C���m�	�)S������>�Q,K�7�n���Ӹ�D���I���^5GjX��*�R,�a��Dd@�B�g#��49���c�T4�~Wf�Х�S˞^�XV�I?U��k= ��_��/��k rb>|��`�d']¥c�ǳim 
Ȝ�_�`m2tcԽ�<�@G)4��%jK~�0�m��g`*�tG-G�<��
m�Q��5�08l	y�3�|G	���d����� F�`��3�KTQ~B}+;oHԚ��L\�!p�S;p�Aqg�HAj�@^�U-�$�oc����;��`�"�6.	�4�|��C��n�a��[`讎�2����u�,U������ȭ�d�!n]�&W�,u��)$�a���bk-5k�@����ԧ�?�NӠWA�HeP?f��Z~V�;�(��:��5������|�a�����������O�Ǎ���f���:H'�ge�\H(�V&�[�0"|}pC��Q����P\{Q�ńP��JurЁ���)#3��m���i�R(�
��H��uo
�}�C�DXgH��=;1��h�t0�{ۍ�9P�y� :3�#Z���L;���3��*������^<�����"����J�P+cDy��,��R���3ۅ,g>��~	�pmlcr7������rٱE�W3_��I���_u��;U���*B��g@��M*�5����}�w���O�h�[������x+ p�Ao��{&����c�|� /�
�:�c��U���'��P~ ��Gg_Z��X�6ǻ��]'��Z.��m�#�R�,�ABF�Z�i��_�2ǩ� X��Yٙ�����3�gO��J�t��ʹ�&�����t�Ϸ��2�cgi��I�kP帣"��	�pM��(W�[*$�����Tx�Y�����*3��(h��<5֎�e���z���S���Z���RȜ���z�*I|5kH �Z�MmVg�AL ��byA�C�S�����@�`��9��C�S��[Gv�nJ���>�q�n|�v�����>g��h$��;K�En�=���MX_G�]Ȏ�����,0o�/��i�J�9i��p�d�K< ���N��������.O��+��&*��*貗���OQ,��R"Z*$o����o��i�XO�?]�z��AFYSUMXb�A_����>,���\z�i4�Sյ� ��տӇ�w��O��Ur}��l�Lp11�Ez�v+x@
�l�ia�K�}�-��N���"bG����LɎ��_Pý�B�(�B�d�gG��eӣ);�(#>FW��Z�J2H�d����?}�v�����c�h�gR��8gշ���1)8f"޺F��4���Kwh_4�Ô	�jm����a�5H�8dދ�Z�O���S����^����JA�*�{8ť*/'0Rd�A�����XJ��,��_1Z=ஃ�K���/ｃSUY�z�&o�:��%���D>�xr��eѸ��n�]%߼�l��҄	(�o��v���|[�fì�uG�Ͻ��0z�𣴻�S:�y��͊��z:s���������׵�	�6Ր���~�g`�:M�Y�
�<�hR�q̌܈��q}��d[��}b,/�g�{rX�)s��/�͐є��#�{5����N�3J��R(��y��2�������\g��z�c�*�.��Ԥ�kI�9tyB��g���͍�I���]�v����H 9����	5*]�r X���晛�Z/��e(��#��l8�ᣥ	$������c�b���>֝���)D��)�^�*�:r�ΝQA�_:��Zܺ�/�}ȼ���=�߅��q��AGN^�w�P(��0�&����xF)9�ϟ�����~ S�L�X�>�q�j�KJ�n6��
��a��n"IV���]NQ2��<+�<�Wm�&m���U�E&B�8��(�B	���Cu]v���`��w�D��f�]�J�� �)"�	}��8 dw<}±@�D@�GVï~��e��6g���R"�i�Ew�/ç���v�%�0j��qƷl�C�l��y]� h�"�-:i��/E*�Fo�h�A9�-�3as={�m.噣�
7�C��6-������(��Ƒ�B%�6<���b��4�;�0��?3��B-]��B�(ݠ��2(yE��Xp�,u2�-��t�/�>jb�m&urBޫrX�;磱,��H[R�j4��@�|n��Ex�9�a�\Ը�����B�EI-����uWK?O����'m��L���F�G�=~d���r�4�j�0���̓q��6����W�>5'��
I�U-�q��	V�..�`(8n�!)\2��Ȋk��M��nQ��b�@Y�67�0�`�D�О�=ygd�S�J��b<����A�^F��8�_k#W})t����,,@�Q�	O������},���B�O�vv�X�C�v5Z��½|�, �!E���t+����$c��F�FK$�3�����]S�>]�M��D�����*q&Wh��u�?���Z���$��
YJ3�V߾`�R��$m���a옍�>1y�n�m�L���-/M����#x���w��vp�Kp�`��V涬�ީ>�����u�5*�$*�W�(>P�60k�m)�+���H(1���k��(��CEH�O0�n��ż���SԴ͛�����&ć��9�q����rH�0v_�K'J���$��s7~�R�'���>ɀ�}�K#�S��ͬ��7e˖��8�9�GrT0M#h�M-{��+9m��Ga��k��l2��I�ms����;������J�OZ�Q ]����U�k�������O���+b�])�m���� �����Ѹ�Ω���(���[��F�4=c����k��1�'Z�Tm}��Y�P�mf\_
a�:�hK^0�J
bO_�|��G�E򬺷�0C���>�+�)c�a%�.V��鳸��K[0yc�LiX���	��y�;�CATe����9&;�H�������붌Lz�0��T&�K	(�����h�;c�̰L�����18!���<zꀰ}\#lk�NY����T��)o;�Vbrh���(���ѧZ����n��Q���F���gx�[/�MH�z�X������~��^T�i��b�����OC ��f��<n�3A]T��\���?Q	T���9'}?�w"x�>TK���Shb��A���ůp���zڔ�t�La�"d+�9u��:O�����(H�o+ x���G�rǛN�J��t���̭���dt}�9'}�c��y��&Ⲕ@ 1ő��Jxc@�4�X���3���]�#�OfU忞�"��'��O�뉜׮�.�"i�k�WW��5�6���������U�F3�u�[�I�.@ sV��HËѤ���66X��{Ftڃ�@�@��&X[�	�V�J���y*C��X�ShM���w��K��>��$>�dpו�xr�Ի�oy�%z���6��ϯ��$�:�����҈ȟe���&D+x�#��\���a`� ��%imQ_HԈP�HVS�������7�i}#�r�K2�%qψ1��'�+�9S{�H�0�j���=t��#^\�T3�ɓٜl�:��pʔwb�;F�<� *R[.+��Fؕ�`'y��|5�dY%MZ�l�f������DN��O�)kR�|.1�qb�T��>.�YwEz�����Wi���U^C1�,7�����L}q���H�K��5��2�p͐@B��S�_M�wc �Q��[���eM7�$��1"�h�c�C-�
�M|�)~�F�"̀��)A��uϿ^q�s݆���6(&�x��? ��;!����FgEMۃQ�X�D�l�mdH��VU|2�f?����W��P�1%��]�R��xu a�.(���������?*�S�[�s�^����*��81m��y�;��󠟳��y�$�x��x�� 1��*���!��lCZ�_��#z��Wp�F'�iRi�9�싶5�aٛ�W){��W����ᒝ��\��[MUb�Wʳ�Hh�%����Ou��y\;.Z>͕����$筨���6���<��׍@Yv�I�E|�@@{�;<�ѥ�A�t��<������_q�;4�����?���0g��3&p�|"cm�*�.�����f�n�;�r�L莂���������N�c:7g�cVZd��<�ABjez&?�ӚӰn����ǼE^�{$D�L*9N�&��m����w�]�Ӆ�֓����MP��b���t�<C���U�(�UG�`�_��X*�]Ct���>� �$��C,��d��o��m��h=@W����`_h�+�JO�-|���*�\|5�_�_��Z<喿ိhs�B�QI��:��bk�_��=REϔc+8�5����P+'����I�-K���%S!��ehug���m����A�)7[_#��Q�����Y�
���4����l�B=�������N�����ݟNR@���6���\%k�Abm��r%kT��q�6��x��o!G8����Fv�_�(�I�~��X�#���ƻ���7Nq���C��ɩi:ԅ�'8�z��\�Ĵm/]�7��Sn�g��' �zTQ��t*��gN����ހ�����I�K�IkE����-.�b�3m�R ��=�<fc��_9 �u��"��)���:��\r��IO(�͗#Ϊf��]쌑�����'J��$���v��Gj57��%0����qV/s��eE��u�[zD@?��;�p��Ƕe�I�§�������cqY�O{��{N������64�{v!�I����H�#]>+}���;g�@r\d�l\��R��4{G�42*#9�q�
L�����SFI�(�B�t�=o�]��#�"��;�z���q�$m�� V,��gbѲw�;�b�+�[�]�Y�Hp��|��`h{a�CKYp.>W%�"�(���7��LЃ�y�H<y��(^�&�VF���0D$/3ξ���>!f��	�XZL��x:�J��G��'QDޜ�7���^�?sv�sPƂ_욄;�ܙ�p�2�4��e#���h�`�����~p+��(�(V�9��ˬJU�˂Y|�!&'8ZAA�7Ӷ�K���c�������O?��m�}���mm4���eJ}קƶ4���l�Y�u����ԙ�:@�f*9^������ߗmَ 7�e��⎪�{�#y�{g!u]
GQ�CzM�%)y˦�ݥh��]|�i��㈮��O����|���Z�	����_J�;����c5*Ǵ�U%�{������N掄�&[��զ"dȐu�lW��Y����5��$o���h���v<c����τ8"K��$��;Y�����j����;f4O;�j���t�R�		�r]��F�$���J�:,D��lm1�������&i�S6�(��-O�zHN+�:��q��뤇�k���{�q�Xk��f���6+c�}\�1��I@I�T=0��-+��φ}�}o�jc�YW��L��%;Z�y/��5Α��ӯc�&�Ӗ4u��]�:�co^#�_W�b�?��}�`�A������x���F:�}�ىvpF��^|ܒ�[`j�<�2oA�����[s��g+�Փ���A����k&�D���/7��+i����J\��hy�*��*떌rD�[��w��M�5��
.��R�J���=�lQ�z�ăq��0��0N����-ׇ@�+ou��8����ԗ��������=���}����Ϳ��^P�9�	���g|�8���5<��h��>AQZ_�쮞����,��N4��Q��D+�q�Ҏ��Gi��,7,�/�a�6�?0�LO�HO� 8������K=CG!�5���2)L_�-dU��c:�������B��@�ǃ����Dr��+���zg"�JC�xF-E����v�|��y�`ޙ�HafR��tY,8L��*�zTAm�^@xr̎"����M!P)��	��y�.�=ڑ �z[�;G�E�{�ݙ%gRy,cr3~O�:�
����C�ٌ��pл�
T��z���(Y{�_�ô�4��&�YOw�e.��M?�	��9ʰ?m Jf��G{�J���g㵹��}`�Ik�#�2﹡9�O�i��:E��3e*�j5f`9������a��/�n�A&�^�ǅ5�E:�K�4��ѥ{w>bb.ML���0��e�eYz<>Sk:Į��x��b(���ZI��K��I�xڞuh�5b[?+��؏����Tmo���a�=e4��d�x��^�&��}���Rw�\���ξ���79u�Ї�X;!&��ًV\T�n��e�ηF�2��3aK0X�g�����ʆ�d��@�Q]�Jv�?���q�Ξg�mB��n;Q�;�c_:�W$�0�Ղ�s�;NW��U���t�����;Nuߔb{�cw�ځq+bDb�ۄ`�젱X��:���,X���@%���4P;y74x�71=�ߑ��G��[�d�&���Df��`jFW~����[\��I�׷z�b�0g�v8C��'W�=r׌����%KZ��5�<h�r��;D��e��ӱ���'�-J�9�w�^����[̉ ������0�m̓5N&~��*�������zߞج��ԚOO�\�M�_- ���qJ�d�ض��;&���t-���\xf�c h�;ߙc��Y�BAd�����uy��Z��?���Ȓ��d�f�/�%9�]��j!@��9����h5l�E���L��Ng�l�^�0����_�_e�3��Q'ϑ @I��1���x���2�R��s��@|�(�
_|*M�G��t��#F�@��c��:�C�}��`՞5��16<U��֞S����7g��w3��>���/+����]�+��e�L�d`�I8�z��B7�h�0=����8uym�ق�4���ӻ�����X��f�ќ�sٶ��%*���~��}/n�����>���+X����3M�� ��� �V��Ɣl�b��7��<�G�e�a����d��;<^Js^�W��x)j����Z�� &3���qKn�ӧ|�����}��(fP�I��?gr}��kzJ�!ƔY��ݔ'&���UN�
��z
�\m��[xxŹ�D6�&^�Y�$��t�R8�8yԖ �0<>Sߣ6�?����K�ߠp��?
;����~��hn��b��s	�*ynW��ʦ;Y��1�e��c�G2��������A��7to��v���-��u���YCi��{;��ԧ��S��\i�A����d _�C��z%v&�ȍ-0g���'5 t0��S�Ee�<ߪM�B���/����3d�5�7�ڷ�tI���owe�<���~�D��h�S�=6'2�4+��峩��2��M5��c���Z�:��+�B���VK��Řk�*��yi� !V��`).eRܼ��6����c�Vg
h
~��'4.�WÊ]�]�sy�xǬ�3'"F�a!�[�m�|	-^IXѭ�ߩeL:�=�pq�o�;X��!=�?yk6��Q^�bFh�.�#���p+l�d^�4X$Ț)���~��u$��sz���r�o�����h�Q�D�)K��`�K���U��l4��u�����$��
�^�( o�4�n!��-�����5�Պ6̟�KWFf�1_��۠�50H�q&(�?�.G��,&v����1�q}������8\�_�������_��<WT�`�ǌ3�_g��h�_��*@@!:���Sޫ���0}���1�Ln����H��L����Vp�D��A�G2����لK���8�
����\	�]�_
e���+bʦ[w��ߙ�8\פq0zײT��6w�$O{��sb;���̌��Ɨڄ��M`�u�oU� OY�&�ld�Q�&/8�-��ԏU�O$�\!龀}󚽇b��i<B�B��]�ButN�!�Ӛ�Յ~�w�%$<ݥ8 &ݖ|k�������r���Q9kA��W�k��)f0vH0��&�Ӷ3�IT�����e�t �6�p�˫Px-������:QC�#`6��S����>��k�8"5a(rz�LH�s$D��5<����\�#�S���ix]�|�{�y>0q'���L��*{�Kwm������J���)�?��5���r�I|wv� %	Z=5��o�3G�l��1c���\Y���}��"A��!���˰�P� ���}�͙�W�갉0�8kM9J����ӽ���eP�T,K��jWnG2s��k���AI-�V��jP+�M�b4�Y��&�oF�e��0e��+XLPcq`�H=�_TS��إGq+�@_��%�rK����V���^eJ�g���Y_|��.X������1ܒLL	�2��4����*U?��K���A�ߙ��ș/��$C)5��W�kp�c�kT��S�TęV\QgBeQ��B� �E�=��Ɩ����F<&�-e$>����W3�n�Ī�PnW>�zJ7ny���-S���Ҹ�2n�G[�"#O���L���`�6n
ˢ}ٓN�tP��3�@;b[W��H����ܞ/"'����&�B�$�wľ���*g�Z�wJ�3��|p�۾��@�u�ï���#0�Sj+%�EWk�4�GȄ�0��C�*8�K���O}�1<VC�X��ɧS�p�*/84��cD�/�{h��d1e
��x-�[IƋ7���S�$+C���s��q���e�m+�$�h�Ӟ�o�-�>;a�QeUI���H*���(��b]���9[N�ˡu�긼�h���.�"�����8�� ��ɯ���վ�H�k�DV�*d%J��K�D�O��c�V�X��<U fq�\G)�Ã���s�jӤ��x�ݛ�jQ�����K���:�v�K0%�P�5S�� _j��3�s��S$�m�(�:E��mz�&,�cF.��2�6J���+���E���d����G�w���PO���jL�����B�~>6Ѭ$W����8\�*���>y�����#��!�ɚ�!�m�+�Q�xK�'�5=�5�"t�e��E&��_�d��:Vo�6��Q���P��O��B<��>��H�pX0d��y��Yi�윗
����3�,0�Ŝz33^P�t[0cm��a��r���r��i�
��LSF�U�N�([�c}I�zr�#��sd��#IuN�_�f�$�\��;��"��g^tb�5ą�a�AB?U����ƴ��UiuA����0C�Hrg��n϶���<�+��%z<גl����S)��$�y��-\�d!����w`K���%���I�
E�5�C%�䗋q��|�A~�Y��»�f�r�&
���
�]�6�]ѿ��]����de���`��f�ko#��R?���8}{�?�)��'41Mc��q�M�5�Y�lG�JV���d����~f��r�DV	�i�OO�yBc����B�Y�\��g\	V��=ϑuQ1a��*�jѵ\�6���tn�|'�S~!�>qX}�*R�ʰ��؝��_9�%�Tw�`g��9^Oni��<y����P���/��Ǯ�2����6s��8Q��u���3����6���۟�6y�����u(�J�Մ|}��X+B?R�mn��cë�:�����N��b�iU7��X��|N�����_@�]����z�e��+d�`�>�ǩ�"�l�OOcN��VB���Fe�c5\&Ё����P��;og�mZ�"0&�qAk�!d�=���%�n\�&�6t�c\�y(��Cf~�􄣸&�����o�7��jWY���It�/@����eDV�I7��շk�\�+��a �U p�ךH�?DH�>���}#^�8�T�l� d� x�U
ʔC���D���E.��~M��4+uE�������i�B3�d�]��:?r�]�Dy�o����%ԓN���{6|˃5��d{?�a�������?��1���o��2��x�jߘ�ɺ��Iʺ}����p!XE�������6����9�)����L�m���x`�]�02�8&��Ė�Eu��>�˓������fn��L}c�(�Z)�v,���߄b������5ld�!���ǟ�`����zL�ce)l;����>�p�	�/�^�^,�O�_~�y=��E�������[^�׻�Ӧd��6�E"^��_� ��$���m"�(v���O
��ɅF��?Nh����x̭2=ŗ w��GT�ش,!������q^{��)�����'{������V
�����s��]���}X�C� v�t�cN����F��E�k�5b5�}���#`0i�)s�En�lB����Q$ś��Ś�yٺh�{i�'�֚-���ˢ辯�b��^c�X��9��i�`�l���.#��4Ǎ�5m�΃�}�T9ڽbnjP_�t �+��_6Y��!p����jE��֜
)?�"TX��<�{�y��)u+�Wl#q(� ��!va@0�}�{k�e�|'c�j{��ts�u�b2���ť��J��.��4/�E]+4��6	mM�������H�(^B���i��3���X��#�QF�}7�;"��f���t�j�=xU�h"��e%-�lp��ʎ<���ڞ3�)f���>vc젙�>(�v��1��U@ĕ���m�}<)k�_�C ��C`fC#��/�kb����C7��Q��b�?$���P4C��0�L��XEd%��B����������j�n3�
ցOi��H����g�0������fs��gQ��?Y�|������T[�(u��|Q=s��X�O7 �dN�ۂz���������2Y�ӭvՍ��ǜ�+@^ת����:��@ۀ�EG�]۞"�¡	�mW��Y�ⶻ(x�P����,�����B'�3����I�~���J&i�������O�"�����L���"P=-��y6�p�-U��(�l�? ��i1�5m?�c���Ռeۄ������7�>%��6��+���k%���˒���A�(���/9<Kzo�u�&[k��!{O������+Ը�Q5Ò}���T��5�yW��oĢ59m���F�2A5J�OK�_��n�B����Ǫm[Z1����ą#�<��F#)���w���~�WŅe5���ܣ?D�ԩAʻ��L�2�����m�1�SK3�XJ�x�.�)�|�,�Rwn}'�AݓU��j��#������1$�)4e/�b�B���P��0F.��@���XG/��n~α��X�@���laū�۞���g�b������F�J��.X?'r��i_A��jق��Bz�"���q#%�P���������E
�{��$�;*1�W��W�9X�X1n�������Y�*Ǘ&�XfE0Brh�;K�1מ��e�/,%�l*��$�~����"ܐ�`Rg[��,K8�]���P� V�����
Of���Bj�5p3
���7R���,׫���`��l=�P?{\����b��Q��琍��x3]T�@���tPᄉ�J{��l<���v���"�.��b�:lf�y�J� )��N��<BH~�y��9�w�k�+?na[;�J�D ϼ���>#)F�v	z��ѯ�*�u�������$�o`���Q�K���v�N�Ӻ����}|:�?�M3c�&#\A�;(���4/�1��uyV�~��X�L�>� ζ��2��$V|����x�>D!%���%���T<�婣v��R�(u�Hc؅�5Ьa��	�*J����J����b�F�\T�2J�L� `q#(� �����f΢�0j�"�O�)��>��>:�����r��.�T�!�
l8h���8�5��'�� �E�^V1�ѯ��eI�)�1T�K���
�<�̕�.qu&�~�S�V�op9&������߯/��h,Y���E�0�WW�)V=&���e�0X�m���Y2���THEy������V-ܞ=�ǘ�G�2�}�@���D�,̔��wTL�����M ru���ސ�LC\�UfQ��yQ;�D��.�)�D�z��Sҋ�/�h���������R�ݵ�`A���@4��ɟ 8ED��35�;Ƽi-2\����mz���Z6ḫ�=��ϐ��	o����V=߂��P�P�+͆6��&��_`�YV�V>��X-��M��|�x#+���`&g�����bk�N���1C��A�7`}����N��U��x�����s��>�*�����'k���ԫ�O�%� |-����bE��_Ik�C�z�s���C�H8�h��6��c�8�cQ���+g�O)�e�.`_�砪��?C��LvbԦ��1��^��KOQ/�� 2�)rj��B	ǘR?���79w���d��AhG��]�;��8�a�l�Z����t����RÑ c�pg)S3`.EN��qE�<v@��@����)���%��z����A��k�D��)�˟�����@H�(�w��q]36�_d�ǋ�N����w�\�{7p�/�ήC�ɭ���}Ƌ���ac�T ,�7�ˁXsa��N���Z6��xf- Dw&Jo�1!��bC}��i&}5%��F߫oWM��Wm�=����+�쨺���`���i��C����v�E��E�Jhs�u<�������Ɛ��ґB�9��xE�����0��S�׊�r�!����x\`r�������ŗvAe'm\Dݘ���hje0Q�r�P���Ơˢ*1��{�({pS�˖�=�Xs�
mŵܳŐ���h�'Ԝlԃ����-`̧R� 	�����	�'-�/��c�N��.�b��"��ņ��i7y*�"��~]�%��۾���htA��[MY[P�6�3V�-h_�Z�/B�Y@���S�zF^Ў>���	�����3�ٍ_XߜQ����	,�HR֏��|>\'	)��ع�Um%S��P"nM?�b;�kpo�v~2���iV��罹����0L�b�=ʛӵ/���\t�|�hw�XÁ8��zjw|��H;X%KӅej���v�	�����Pm,a��YP�r.y�$?��
I0h}C��.��??1���ތ�S�D�����A�/ts����Q-3��څ㵥��Z�TUgJ(|��⫄��r��8�)�U-�� CՏ��|�Gx��ˊöWYqS���s�rLY;2�cH4z�W�����aq��ֻ��D��"G�O��	1�y����qoRIMZM�����	�����.��� �:/3䢬Wr���Qci`2!Ig2
<���=���ُ���Vo�XSn�P��G�09w��i�lt=l��^���]�B�wg����Y+�Z,h���J:[�}M�vs^(�ZR��|Hf�C'/Nq�\��4������rSr+�͠�>]�p�)>��!*{��c����1)�`�v%�F�ﳔ�9�˄_��n�a��b�����:�U�@+��*XT����b�h�to~B��ߒt�,����z��{�<� D��>s0A�q�s��&���"�r�7u51���3˖����A�@V�]���U��@z�o�NWO��m�=9�H�h�h�@����ffZՆ��
�@��K�W�w����~H��"�+E�g���[S@3\�j�RD��Ur���%��j
�c;k%�#�]j�y��R���`'`W �}Y��(�Y����8I����ͦH��]R�w.��րAǆ"�ä3��΃�W�C�/�ܓi�j���X츾]����ՠ��O44�L!oO�c9�~r���D`�j�/�skSGb4���e��ƱO�Z#�7l|�?o�����ufH
��Cq>��B�D�@�N�rx�O�ӌ_d�q	��|{��{T�3�A�$R�H`%a���r�G�%4�c�xo���q�r�c3����^�������?��5QLȾ`յu�o�`��N�����@�-��4J�Jk6�jѝ�E��H�
ɮs�s��C*)�a�,A�piL�DR��x{�����"g�c�v��23`-��t���X����_�׍��>Қ�2���^3x?:�_{�g+�j:BG��I'E�B��翫ksŗ�g��g���I�lYGT<x�yg���r�MDB��mN��igst�2�������4Df�)7�h�¶А��ꑟ�\��L��rp]�x[-$��b0Ґa����@T鯘��ۺ�-�s&��$��P/ñ�o��`�[8��S�{֢r��el��F��ĥ̓2-=�%9�Z�����h�����7��3z�nτ-DS#�/YԐ75i�����`_�}W�y���QB,6�Z�2�L.<�߹ڰ����+T�g���#p� �� 3�f����+IH{��S�{�xG)��ᵻS"w��Lb&�ô;Q��FD��4=�� WY���3��g,h�.��1��ꮰY"�4�\"̀td�u�4��X�O+U@$�OGa.�.R[ ��g�Oؙe������-Lc�]��P�dQ�ͪ **�����C���DݒA��_w�#2�|7)��D�,� qQ�Q���8�H����P=0g#�o�G�\�:<�܋�L��/�#�%��P�gq	����\N����g
�2T^䏓��i��N�xws,t� 2
�;��a\�vc����uO�By�F&�I�q(F�]Z�nW�l"v��\|;��e��Ҩ���T. $(%b3����X�r�Уn�Ot�<"�����[:��(^1z/�Ϫ������W�wDM�o]qӬ%,�UDj�\�)���Nx���8Р�Έ6���T����1*I�GD�\R��&e��)4j�����\�UX����a�\�E�>����#��;ņ�n"��n��l��NPߚ�ϖ���˝�f��ΰzƲ|>o ��"ŏbm3I�Q4-c�M�RC�]�� v�,�a�I�'[m�*Ҡ�����7c[m	+}=�$Ty�Mo(s�d�����A�q�$l�u�9��TD�*Q��m'��~��L�%�m,��#	0�D�9�-B���'S��:H.-��.���f�_/�J���(���_7yjE��AoIf}�
i�eX�"��PC��7-�ޡ�K��:��V��C����ƙR�+�iw�,�"#*�ψ�otA��Vo�ƫM)u�9�R7�j_�9lO�~�As��Hh�X6� `�����c������^����cU�������C��6�~����&�w������ Ț1��T�?27E�}�q'�];��O�vJ��A�� �u�q��䟨�|K�7�J!���)�����������[v����v3-)�[�%��^����c��oQ�����:��Wa�Mc,Պv��{��K�L|� W�G`|���Ð w1!�ά�p�J� }��+�n�SL�p� �:d(4.��E�lB�	[�e�q��p�S�%&��kk�������Zi{��/o�~L,�l{ K��|y.�5�o��8Ï�C�8�)CU��0<��o��]�A�Y��)0�b��������%I���ndz��������е�d����X:"�
��3�����(�S�?��,b�l{��_�z�!������E�p�|�M��aN�	̦NbY�;0^�ZCvq	HXsqm��}I#�l6�,e��R���ֹd����4	t��9�q݁�]b�J�=W��s��I�(kNw	�_6l �l��|�2�e����)��,_�[�(��T�fi��c���<.����K|��!�%�B]�vG�2c�b�v�� w&�i�O�]et��R�nݕT�fJ�A��T&��I���q68�!0�f��.n|��z�-3aS$��?�5�ծ��
���F<�����fdb�B�MT�����uw�7w"=�vg�hFq���$ә���Ce���˝��3F��z�j�ضN`O��:�n�o.Rh ��}�����i�����z1�?m?��-4>�����������o��D�����)�4�+<I����ANw��2�0|��i:�5
M�Ϛ��୺h�ʩ�V0p�$�uŗw$RO������U$r^���:a-�B����[Ŕ�P�������E�#��bC�]�����H-�
D�Ӻ�CW�p����W ��oh���Q	�4R*3Qk�*j��b9G�J�H-�S*D��~W�����ЍU?q<Q�bGZ],��3�WF�Z�.v`�t�D�<_�oem}[��u��@�?q��1+�������`<*��O��'s��h�]���ʏ#ɦ�M�DwSr���
<�~E���h������UӲ9��'�����bC5#^=a=��
J9CK[d�Y �C�f������������?3Ԉ>}v����4>�����<��J�`W����j�.��_��&H���6T�$�b?����vZ�~�i����$CJ$e9��I���\d��
�T�b����&�`��P�[w�7�Ǳ��c�g�(&�{�l�7���C�pe��M'B�OIb���ʻ�6"�l?�oɌ���4��M��Ւ���rrpy ��l�;���Ǳ����Se��>��&�����^V���l�����pc(!~v����=<��^P���N�	���60�����*��EU�<�s%3��^;�^��c4&=>k��1z����Q!�4:�NUhQC�i��ٯe�}d��Ei��X!"3�h��2'29�g�-2�6x�ם��$I_R}������bkl��z��sP�V�U�p�b�-Vv�&��	Uz#;/2&J���O�i,8O�w�L�m|M�V�7v�ksRJ�J��bĔI�{*���{�?��6������01�Z��Hh����O�q�����GTڇ����^�]%ި�%5WX&�AM��&�b�)�Ğwp��奃O����%i,�b&m�������`��d1��'�}�Q�e!�h�$���σ�UE��}���n�//6�AR�ޕ��ˤ�N��+����X���『j~V��{h闀�9�x���_f�'�׾��J�ʞ�&�����]+�K�1�D0�g�Eļ���
i��9%u ����E��S��3�
,&Jg���FR��c4�O:$ȸ%�߰�)��8�V3Oϧ� ��.�6J�Gp#����K�^�1s
����%z�5Hx5��1c��-08~�E��ߤ��&�Ɛ��>M�׷^�S@A�z�a,>��#��v�	���+�8 ��G��,Ao���)X�N�4������0���`��;�"E���D��6T��!�B�hV"�:4twQN�{oE���>n;l��x*�Uj�U�OG�J�81�C\�x��P�n�B�|l ���ؑ�a
9�N���@ �J,��煶��L�?�"�g�����Q)��cudK���
+Xp����:P��OqS��M@�J���ߥ����Ie\U�b�-\��Zt�vݘ)�8��	R�$�P'*O��R�}_���s��8�e�M�2��xUP��;L�J_D{Լ�n������mܕ*��W�>q���߾豐�CC4Mn6��+�
�$��ͺßP��Wę֣K[��1��.5Ѓ��+�����`��,�
��>��r�Ur�DӠ��ͱsY�QXw0C���,%�خ��G@*o"��������t�|��\��,z�;<~!e�s���GW�m�_�=��J`�v�O a!���x� �o���Q�
&!(�(P�s���rtA�gʚ�xS���/ď��.N8ݽ�n��U���`i�����	H�}�@By�6���Ⱦ}���.�X�DNDۦ�	��F99"���&Or��Ҿ1�_�����аB,*�.�G�X�K_ܡxO��?�B��}�ۻ8�vvF�4��OR���%q�X�H���g�ON���i���q���3S�{z�}� �bja��eN<����j(��z'1".`S��S楢�q���I<U9e������E@c��,�l��u;L0���z��|��*N��c"��]����YL��ӣS2BbPz^�7�(����Xr��g�@�N=�A���䟌�Y6��8d�� ��"*QL9��k��^y���_ 8��D'� �m�M���28,�i]���Qr��R����D�쯯��(W%7t;�6-������K����R�ǲ��{oK�l.}�ѡ*�r6@O߯fCK�����w8�����0ӱ��i�W��F��ak"x��.��8?��G5G8�1��Ymy��G�,���*�V����2|L�sP��AT8�o�'2l����5��Ž��D=�c���j-wR���9[��%���X�-ﭭ�#����C9�%��b���X\
���OcxM��S8���0FkW���E����������ed��ߨ]��?Y\xG�EȖ釹���w��+<�l����6�(�����K�+q>L�1����O�)2ϩ4�:��*�X�hl>0�:��V;�l�����Vt��Tw��Q�$'ٓDX�\z�� T��)��A��1c�3Q=�:K[�%�H���i��?���?I���<LTlߒ0��vUB�Rjӣ�A���>֮a������@���v���@8�|��U5�%
�I�*�!WQ��A�T�£ۨ�<�].�G��hW��\-�P&E�IF�n�w��gg�V22���s
_��\�Ka7|�)�<P�O��/)(d��xfg�;��ʌw�}cX�'���i�F���D$*���R�ט
I���pu�K6]G�A��0b64����1��#��\�d��c�F������RD�)KDx��1<����q�ߕ��D����cx'�9y����C��.;�2N�g<K���L*��D�l[k�;�L����O\">Ց�Q�s�]?V2����<~�6`��֮%ޒ�����k�`\lu����d�k��e��@A���;�]X�mx��� K��]��T�G�&49J"$��2|�m�%��d�i6�н�_�{���ɔ�������JR�t�t,��B?�UEߦ�}�J
�Nަ|OX���Ǣ�	b��?o��\�F7�d��A�g�+�ng����Aܓ� k�������y4�X-�J��Qt���>��n�HJG���������p�I.|�J�֘D���9@�V�����;���u����[��&/#,/hW�����h{�p��� k����?aU�џ�q�gi;s~����H~ji�r|�~�n`��-�^�����������w���gd�H-禣@"4���n���'�R��{ײgl�>a�UzN�yt6�(#&တ�X :����� �OPӄ� pK�9�MX��p^(�iG�{3��d��̶DQ�ME#C�Ҽ�����]O�9⓭��\�.��$��`��G�G�)�s�ɖ�+C�"9�nN������_���5Dd��,�����B׫'�EU�v[2-�@�u�k�\�l� +w	ioX`�&�������xU���q��&�����:��
���A�鄦�G�iO��5ނq��������"�W�I߃{@G���)��_0���%��1"�7��ږ�B���׆�m�>O�{~��Ù�9k_���2�מ�?�k�U�m�~X$�����@(Q GLy;%|k�S���x��9�-�n��C�PLw:�in�gpPe�װ���Kn����4�b5�J��0	��KO�Xa#�y���p,N�[�M��'�2�3B��8���*�����_�k�y[�����eI��Pv�l��"��/x o�V�9�nr��=G@f'Km1r1���/�n8�@
T��� rK�ܗo�V������kz�evRх�"�PX�Pf���y}�ٔ	a7s��P@�S�Ō˩��XR��l��sǎ�$����i�șS�X{-���l�A {�NN/(o�y�ݧ>��ǜ�	?�bR����1���n7S�=�ǃ��5;��6?4+��f"��I[��#�Ȃ���
��(Ni(�4u�Ǭ<dOߕ{+xo@nNX�C�T@y��^�!e�l�D[�X�c��P�t��^��W�����VH�ߓ_��C����_��+�8ri��[��"	�|�0f��J���߻���6
Z�� ��>�N���5�U�����뫔�,[J~X�%�_����-������(��FM��gZ~Ԟ��ϥp~ <Fw7#�JGu�k⮞暻�#}������]M��p$���A'x��;������B��Z�TR�AX�^)7d���Re���uR1���ate2����n%{_x�ċ#'Mz��-�����qy(k`��02��l'L���O�^s[���9A
pU���t����/�R��������!�"r�~c����~��r��b����%G�y/@f����l8�yH�� l�ڻr���m���Ti��!$TW� ��
�����	v`�(	_��n�(PA����j724.������P��W$��_� �v�-g���S!_�>Z܊���7/�i�+��v{a���b'�8��x�Z��1���}=��t��J�3���	�����#�s��+|/���1��S�j�
�'���*#�OW����
|��=!l�0�U�.�Y���˖�*���2��!�i����jMBή���r��	��N�2�^�o鷷S7:ԵT�(��By�Y�;m��PdΚk��R���Qi��,{�����Ex.�a� ����tCÕ	��ș���^�\܆�]?:����m~�Ԟn��OP�z�K.��DOVm��梍pX���rd�������
�
�?t*�+���]z��|ӿ,��Q�S���aWe?$����~W9�<�|t9�V�g�4yNn�b�����NÄ��	���?7Or1yҌ/��#���c����5��m���~���)���,s�o��Ĕ�3��ϵ	��>��o�[�8�+��W�AA.y7o!n`͒
�����	�v��)gյd�j10M�-(0��Z��l�,��JA�%w�N��ڏ�dnv�FS�C��[���i�Ȥ�㯫]���}xF,�m���_��	��(�fIL)���WQ���s�~�`@����\��3�.n���*az�e~XVm�?����cG���*�����a���W{�4I�f����u��_^���t�]ȖAGxEZ.���#w��4q�B�z�δdX5��n`�O$r��9���+��F}t�������g���.���39����餭���s%�+�X���\|���S�3�LB�j֥�X�N�HQ'�?ʈ�� J�ٓ��!�6��1��ۭe����z�ӟ#�'B�A\1��|@��-�R����D.�(E��������Qr����(�O?�S6.D�d�X.�& '.M���O�P�	�١3�и*i��:���c�����"ʔS@�%��?G�ҟ�L�Xz0V0a�1�r�&�@��:��u�im� �{�����e���@�B�� @��/�>\x�U���f�?�"|��IE�^OF3��<��L&pr����t�t���GUzGbΐ`�ܣ��ى"Y��WM���p�^�N@4�RTU� o�`�K��Bjr����;�k�aҬ�ʿbT�\/�'jҸ�I�'[�Q��zv�/4LwTܗ_���=������1%�'A����\Z�=ě0O��������p` �����EBXQ�a���q�?����z�켄��,�������5����!�rr���gM����fg#|9e7�^>i���nG*e'�&�m7�j�j����X�AN���k;s�R�$;lX�nr�IlS��t��o+�lU�����A��@�g�b8�05��:�%���PԤ��������'���b���K����Эn�~�G{�����<.���a�5p"��I�I�Y³���6���Ǡ�͕���3��H�|7K��PD��Z�U P�XOL�q'�&ٶ���j�g��{�QX���q��<���-����%��1�n���y�
.��v��3�Y�f��'���p���<c�,��,��U���K�%&��1�
�y�p6pe��0\��N���>�1Ј%u.�UX�Gb��>���჋�Z�v9z�7�;t��Jƴ����!�yYL�_K��@�Yq�4?���ļ_�1��'��^��5A{�\�H'�:TvT�����%|��i؇��#�'�b�aY?�XQB����2�s�����-��L�/Vk#N||�X��Vĥ�V�����,vu?�r1S��jwP���%[��i��'�����Ś	�
�݅�a�R)ת�ZJ��PfL>����5<���
��8�Е��l��G.��E���>�G�^��l���M(��)�Ŋ-��!�?��4*���7���'�-XO�Tԯ��vǮL���-�p7x�������Ǜ/Dp�u�'��*��]�,R0��,�B���e^��M; �3겊C����ݡFv�j�I>zV�M�~5��!x,2��`��,q���`E��o<�^!tY�>n:�����8``�dO;jl �1�\�4|[���+U]�����M�ڦ5%F?�\X^2�~�$�#������ċρ�J��ڗc�球�b�K!T)���L�Ϳ7�2��{�㒒�E��e�0hf|ql�B֬y}4�{%4K���z�m��g�a�om�~��^��U��OQe(��ݴcv
���?Q_VP{��CI��ٿ��+�&3��±x�8�!�Kly��;�g�P�@����R���b�k�2 �y�p����OR?*a�W$2�, ř�E�X�R�A�0oD�m��O�$M8K��W�_ت�{L����G�j�Xh9��XI$�M*;�"���JZZh+烸q$k���ϯ`�O���)�~�/��2F	�^p�/8�&⮂���ԸkC �	�e+���m���#��KsTa��9��K3[n���[��0��`a����1O�QHȓ�9�/Mײ1�#}>��6y�G󊴼� �JE��)j�*�y���K��_���7�B-�3��3���i�!�5�=���`ϘDϬG$���'S�e<���0
,�d�a�L8�nJ���88r�_,d�|+u����2)L�&_�{}��WJ���.̋-�z;r�\�F���vv���{T�_Z5t���XŽ�y1�{�rePv�-�ᔀv5.�cRߏ�v�����s�Br7ۙj<��h��k_��i���h�F�=n����7��I|$Ne���ߎ������r�rb�I �n�� V�G�:	Į�~u���6��&!i�G�W�l7����5�c��UM�O�H<8���y��Ne'�6��$.��=z�4��kX�R���rAU�zS���ߦ`�ye}��U�฽�^�QV�+�����{��㪴Vvy��������>#����g�0�]�,��ȟf�4���0>6�K�_h�۳>��v��.(hw�M�#���%U�jነ\&��ɽ��+�[́��:E�j������y寏�|֌y�r�P��B���g4<����:��%,�2���I�sѤ-��Q��������H�m�0/լS��Lf,÷�O�����ǚP�>����D�^�|�6�XVm���c</^^�i�e���{A���?��hb7����9s�����8-|��	9	��|3Ϳ�H�,���'d�+���LD� �����=�k��pG/l�7����#��K|W�	�����ء�(#�{q;d1�Y�GGW�{��	�
�����JF��.2'-A�Wa)\�`���r0R�A�<{�P027�/[�HӜ����;��/�����Z$R�oֵ
�!$��b�]��SGW	[����Lc��$���xƭ�_W_�����[Fix����O��r���[0~��17�?�e�z�"�(u�!����Gk.S�`�����{�'��B*�*R��?Y_Ԓ����$�<��x~���D�oB��=�����gfr/^���e�RÁ����&B���n`�k��AKC����w$��d�a'��CVb2Coԁ�B�(��2�YP~���堵b��*��V����{��&CA���c�3 �V^�12�{Y7%���׹e��sɻ�/��Y�d�|�9��k�Hu"��͔J�����v�S3@���PM������K�9ڨ8!Sp�~�o�q���8�.��B� %�5-�b���@��PBPVY��Wn�1�,���nMpD�.tƒ���J��sۊd�sŌ&������!�0�S;��v��!;;����_t9Aq�:��E���B�Y�׸�g"��oNy�m����R��N�윦g��xÒ!w����
X�]����븄F�~��t�W%��Nq֚%?�M՝d�<4f�N7 u6���/P.5?Ѻn\�D�
���WS��;p�;\�64�Q���.Ileʔ�q܌N��(Ӝ�p�m�E,J��Ν�3�fW=�x��l��<����I�H��t��h�emɣ��"���3��4��~#���j�!�e�śP�<C��7R�����b��dp�Ƹd���?�K���HY��F���lD�N��YvU����a+�?~�a�n|t{��N��`��W�M#��#������%2s�^�2l�p��k�4�����1����!�4>�f\��=d9Tq`Fj9v8�W/��)�;!�n`�,^�"��h|��b�o��B"B�1�c��Ap��ՠ�(]oۑ�%��|H��u�A�/����
F�<����/�C�rP?	��;>�)6O�@}��gk���!37*}�0�e$M������[���j�l�'h�'B�::�U��C�|��[�w�����������m��d�Z:/����.�TʠJa�a�}�YV�n6}����߂]'���M�8�h����OZ�/{E�ʁ����si-{G�|`Q;6�;�?�2B ��~�)���\w����u�nur�j5&�������0p�np0��?R�_h5���&���ъ����.���>�f�l��M�Pl9���8��D�-�]����E���)�E\@Е9�q�Ib��F���C��eبL�R��ܵ܇���;�����_סp����&����g�����%��� ߄iܲ2%�XUp����R[$	������	`�7PDᰙ bߛ�Wo��2
^K���t��O)7bsD�{�Q��Y�}�ȥ�RÜa��eR���VȘM���!4@�(���у�,�Pn�y��כ �Ɵ\�]C�Q� ʓ�4NPF^ۯ���0H$��[����NX�OmRlL�������fW�B@�-�-�_|�I�rf��U�7fȋ�K�(�-�W*� 
|��cɧ�V>M�֨��dK���b��-y��W�-s-|��;��=�nv�eO1$*Eq����2�^����� �I��D�����I�Wp�Î�_���?%605��^���S`2�Hr�n/�p��q�NH7`�La��������դ�D�T~U��T��U�	a��`�E�\bթ�!�������>��O��+2&xC[����eH
�Z�U�	+U*���̛��gҦ��FKP۰?LkM�2�7m����W���"��iw�R�j.��
ҋT��l��<������PYe�Te�9 �u���ɵ� \}x�F>Ω:����rq� �eU�5�E��5c(#�D��Z�,���y�ɼ#M&t0����%�b7���Z�"!9x5N]�Q��3	�"C��������� {@�i�7�w����p�Z������`��u�v%0���2��Þ�xy�'���t��z�����s���s��������xP1���C�È���x׃�fV�HQ�H�nC.]g�y���l����������Gc��dXq�D�HZZ0;�Ds��peZ��Wz�j�o��#����J�_	�c4�n�f᝹�2	M����������i�O�2m��'r;��ʫv�A5Gw��Ԏ4[��<�	+�#/�h���������[ő�m:�s���O]���� C��:�*���+�I�F�Ƅ�As�O����s���`_�a��)�e�L`�@.��V���:G���b��a���u��n�y��F�gZr�J�͆	����Q�>d��fố/�O9mY�ٵ}X�WP��s����
��������/�3�-�ߊ�	��8��~�b�B�?Ϗ-���7�"��y�Z�-�G���?��0�Zx��~��������E������a���K��X;ʲ����a����y�gp:�KjU���������;�#���}����_>�H�?����ċ!���2�����U&� g�7����+��ʁ�9�����<L��ׄ�,�`C�o�÷ �ÅdC�vM�AM�j��}�򇮳g�0Xܱ��W������4<�-p-bܨ�	����)���p��u*���E��;��]H�&�x{�1�;��sk��&�<��fV#w�r�O9���,����a���������i{	xg��Q��2�
��&eP�f�o��z��H�C��G7�知C���$��PJ��ew*�N5o���eBM7��`�%��R��%�^M�p���W9َ���ׇ���%i���7ރ���{��Dn5�UH}_«<T��N#;��W��0AHj�n7ڻf9g>,~e��#�=^�`*�]K��#�א���y��_��F�`X�.��6�i5�	��C�ϓ�&܅�՝��&��s �D�eNVd�����v�*��d�)ŰC�8���.�y�A'$%z*�%��؎��+�8F~:�!��o|���v �,���Q����/̛9,J����gE���P�j溁G\.�v#���&��I�~	�Qؽͤ��M Z��������[p֪����4W�H�-\5{W:�Re���-�,{L2Ҳ4���	��c��50���a�mq�w��a�s��ˉ��?D����Am��H*n�}�"��P�_�}�I�Q�%l��H�p2�1 ����JY�U�b�<v� ه���s��E�f��S��X�=�"H��fl�;�5rg� ������%�#+�qy�Y86x����a"�zUs�UV�|R�񡸖!�q3Y=�bL����<�#�;N6������3ݯ�D�<�zt<Ax	s�K�FCa1��pӎ�)X�I3\�P;�P��uT!�ߔ�2����IP���t�]�|����G �f���|�V�?��Vz�����!��p+�6�@d{F�z��!�a�[�n�4 F}۬3PP�7�2
�iM��%
����{��W6�㩓��2cޮu��}eY�e�߉��0��������c� Q�:�"�Sg�O�vX��9���:7�͚4V���F/4$��.9�׽B��tQ��������L W�g�'�Q$��b�+>K;{���w9jȦ[��1QM�!%�ӈ�	E�V��EH?~�s꣣Cpp�fKb��"�Vm��	�}�K�T�����eK�j�^�"�P��Ҏ�aSA�� �̔����v�6 7�3���iJ��tfgj:j����(����>�SȫH7\�<"�޵�I���䤍��q�12�=SE��}�7ޅ�~�����?2�v;j��^�O+n����Pj���^.�#�\z/�����j^��h�f�A�2�:�_S&%��~v<A��mU"Ո�<E%~�8��^�l],��c�ÑH+ƣ��l0�̀+>]�a�jʱ0#� =����}���u�C�������:_��ns1皲<z�i�z9[˛��e��0�a��B�s����EҚ�zdk_�'�������c���-�������nu���fŘ�.[{���Z]��'�by9�Q1��O�d���K�������8�{��eu��)nՋ��pz|Ϛ��L%2{ �<(Ȁ>@��`?�;QD���'�n��A-/I�����<f�&6�(�g�03��]�f�- �D޵���g<���� ����6m����2�GE�m?�8�-�b,L��mf0g8!���R���eD�*g%7gf�zw��o�IL%�r%Qve��Ce�y�W�\�:�C�zpx���y<B���D��ln�)*�r���:x $�p�ys�J:��+~Ѭ�H=~0NS}[`F�F�0
hƍ( g|�����*�+yu���q��^�^uS��?t�]�er$������g�^�)~m�27N��1�7y��r������&�#��5 ��c�����[�(5��PPg21Z<0-Rn��7�� ���(��j�I�>Pkŏ����e*s�3/,�'8��O�rפ����N���,��>��m�f�C���;)�&*\�U�]樠�=�FO@_A$�101���y\�u�����L֬&l7`ɦ^��b[���4�fdz	�MG�S�#B�����7��/�_�<D* �~4V���&�0#�pW=�C�9,P%��9<#�����դ�ڄ;�����!�\��� ":;���52����-����'1�V�(��<o�D;Uʳ��`^�љW�v$��4���Ӣ�O.T����$ޖI\��2�꿗a/'Q�,[���
�����0�A� �!�a�]�W�MG5��C1(�Ȼ3Mh٦�O���G��їà�*C���H����be�Z�֙���ht��K��W؊'@�+u+K�/'|� [p2���>uO�k�;#�I�m���`�Eܜ����_�LI�wT�al>�\Qn`�jw��+A��@�E<��▰Z�Т��U
E�[�����?����G�+4��!�"�L2t�Ȏ�1��x|��k����xa"�P(�Oѣ�}	\� "c�۲о���aM<8Ux��`������ټ���w�
-�[I>b�"���D~�_�`]��Aw0���})�}e��k��m�K˝?�j��D)g6���Wa�n�@�/���������x�b���ސ��%Gv!��b���d[��kFq=��s�Ć�[ˊ>o�8�H�y�9�E5߫�kf5���N�Z��R����F\�l�c�@hksu��:���� ��]ƨ���{�%i� y�܊��gDq�!�ǽ��oy���@w���%�@ܼ�9YP�[=͹�ݍ�{_^�<�|].Y�����"�J��Q_JP���7��ʿpl=�������}��7�a'相q�Ǻ�$��^-�^V�vi�oí;� �)D�g�z_-x�t�.'_3��?78����q�v��z���r��nS(f1V�B��r���U��?�U��4,�R�a<��ۏ��W�O�{w�n�24�3L�ǣ}�y����0�����\��$��S���|f��,S�F>�S��IM5��L�����"@��Ϙ����}4�_�T�[�3�s�JZ������/��A�4B^�Z��9]G>��,)P�l�z�����N�'A~zv����V"�*�{Pb�� _�ϵ�T�4b���MD����}�3Jq	<n�h�r�s̟~�A$0��ɐ�4V�e?���h}Zu�!�7[�ɢ�о���9��/����j8�K5*�e�ҽг_�����.ғ��u;��L`���{�����x��1��6�NOe߼��qo Z�o;e[�ɐ��Җ�\�1��(k�;�*���S�w~�EζV\��-@�*~�{��yT�e�S(��N��NΗE�]4�;��ǳ����Ծ��N����æƙZ�q[Z��:;m5
c� q�4Wn}'}v �T@0�3�6�DK��v�6A׬�/���u�F&�]������&�T��	S.�:����!����4[��pkW?����P��׻�������պ�d59(!�8�o��9��>��C������-Oz����KUs�!���y	(��7	={=�$���-����TD��]�X��)+�2eu�1�& �I�{�D���=�}g ��U��J7�A��i%*���"����t�_J��U�̀#�L��ļG^��G�=�-�V�L5T���� ���f��m�]�S���Z�g��ϴ3i_�M����N��p7v��΃:9`��jTJ�b{�Ju첓�*xH+@���!;I|�F�Q�6�ޛ�v=�"V��A�N%T�e����I�y3�^3lc��͸|mԍ��q8ѐ-�[��5�l{G��UI�Joٌ���4�����z}"�UW�o�-��˲�s��2����у8K4H)lX�?;�Xϲij��?��o����� `�����9 \��FuY)��%�%�UI� �+v_�#u�� ���*�Rq��a��{x�!Σ� CQ!��D�*K��?�vg�S�q_��1O@-�h�<GA:���[����y�J�|$z%�KJ�@+'R��_%Ս�ꌋ��3�v�\h�\r�xl��(�c�z��u��ޠ#�#,��O��֪����8��.�BCV��Э�H�+����4��am�|8�HG�Xӽ�#3p�#��a�\�>ᔧI7���VIe��/l�LN=X����
�Skg
�wq+B��~���M��9V{��A���@�Z���SC��M�R�	���O��s\i��F�m��z��HyN������ɔ��_�:}�V�3�
h�?o��fvm�Y+�w�����~yO�E�&���tߦ#4}�n�6�3N��.�򈎾8.��u��IR�#w����Ϗ������Aċ(hM\�NP�٣X�A&���)�y�o��A�N���КI�$%]ѴAu����1wr�;���x��T��Ɓ�ʹ��uSU=Y ��m�՝���Z��ߕ��ځnK-k{$���"�U�g�9�(��4�c���V�������F��@P�T�Jxó0��}J���`�4����o��/@5�s�N8ަx��nuz��%&=�P�S�$�{�B+�r"9¡��,�h�ڬ���Ҩ�Km�	�loK
�u�\�NL�uK�3B8���h�%�,o A�r�+�J�9�z��k�$��ة�����F�| w͈ȭ���oA�x�rc�������OO7�.q�͂q��ܮ\�y���p��t%~��]xJ��o�'S�
����0�mo��\�S3�+S����4��(��JZˠ�n�����D��v��)KI*����VWڕ�|Z&���FUZ�n�'+��/M�<px�8� i��G^�����f���P��Yp'���Q6E,:��P�}{q
-������,p��7�@� �Q��OL� ���N�\��ձ��k��Yd����(wS>��sƩ����]�t�;ǂ�oN�� �%�;�o �(Q��z�,6��i~��m�%�~��r�۵��	�3p��h����G�?O�Y��+Y�4c�Se��ٙBr)�R�tB�)���G7�X ��*��;����xz�����V�h�J��h���3a�O�G�/r�F�n3q�7���{®
����C��d���ʿd�[�j�qI��#>B�ү�ZHq��壩� �B��m_ h��Cf���k�mw�����i �A/�o\�/�DV/�A��>��m�d�����;�`^��EO���P��	�)����J��j�Dbӏ�;l�wl�P���v��c�OÍfʃ30&nI����-`����U�Ha��F��'@R�M:-jj�VV�n�2e�0�˰�ƝJ�@<?i!qBP�F՝�'�=� F�P�j�g���.�;�j�C�!��)&dDx�wv���…�����Z��<2q�hے��%un%��o.���u��[��4�e����+9_��PD!��?_��>���.{��S�L��3�����\Η�ˣ�*��apd{{i|�9��H�)���.�cFrO3I�V��V)p����d�K�*'s*0��S��Hm}1z����jc�������W�������\��$\t��a���mˬ[t���Ǝ�蠹iB�(�2?EM�Ʋt�H�'Q�&�_.�4*�Ē����5���ɥ�^5o�t�K���p�p�}>�#�4����ʣU�e�P���%�h�턘S�r��%����Ɔ�s���J��#��e�C5�l$�u	t�zIC��lz��J�?BR�B��Av!R�8�审	�93�Z��?D�~����y� ���E�jj����iɠ�oV���ץOձ>��BH�V'sP���g1���ۼp�gJ����Z4);V�3�T~k�I�m��3^�'�g�}���1�Q�S��2��0����O�˔������%�0(�=�v(Na F`�Rx� �t�������#����+��|�,h֛kZ �l��rA��6O���8�'_��t�� m������K�F#�n���3��`�v�����N��,�IG�j��p9Zn�]�Z�\�[����o��p��߅��_�G�~�'���%=*�4͇C�|v�����X �v��q2ݠ�����.m�/��f6�]�>��\��H>Nc������]X�t9�E{�Y�E~Ig�o0�:T�-_8v�K��vi�L�V��"Vu�����{�B�&v�tgfS�A�x����Dj��:�Ir��ɝ ���,#"�M�@^����X�ܗ��yT���#5Xʉ[�!��q3����_S��=D"�ٓ��JحG�I?���0	��)R�I?�@
\�F��VJ�:���E6�K�$��n|������$�-�E��\�)W�lT�"P:\l��&�B@�D3�-g�DL<8��ch�
lY@�W�vY�_R��@����(i�Yѹ-�����
�%��Ki0#�I����la���&���k�n� ������� ��S}ݔ�i9:��R��6Mƾ�9צ�xZ8*��O���p�u�=m�9�r�L�S�n�e=/zQ1���DA^���Q�Jp7_�ڦ`��'�7:\�o�����<ن�/aa�Q��y�������3�ޒ5&��--���;��f�ax�m+:A3�iu��E>տڛ�!���H�u��g}Пw�����Ow��d-�(ηU҆E�?�U-�P���|���V��~�F������R.m�H�����A.�Tί�TeS���Ku��d�?f$C��[�ӣ��	t<~ϻm��oNSk1��֕-U��%ѦY�Sa�o$Y�HwZ���;��'a���(�D$ާ���I��`��_�H���z�j
1��v�k���5Ųy~�C�;���3eG&����ERPReٓ���(�61�XM&�N��	�W���^Us�:��&$�]4f��ru��l\�j!����D2�
#�م��s8bI��QX�?�  <3/A����O�v,I�!��E�C�[��P�Q�l�+�a����+���НL�7h��H��mL�+���n��86}<laP�R����u�����0��,/,��U	4�����Հ�*�n9=��b|��b2�r!��o*g<�õ�]P�z��R����
�����
�5t�8����x5����$G�o��*�+�s��r�yvN<���̝H��{�E�0�k��3'�JSva���/3��W�D��~EҺγ!�s<�L�.�\A��*3�cب{ͯ�h�"��G�!������nm�k�+�����2Q��OM��Z�b:z��������s3���G"1��f��W�ׯ?.]Ԣ�Ȏ�ct�D��c�<%�:�$af���"��"��ոNp�I�&�}f2C�:�kf?;�eu]Ζ�"�b(1�����c.�v�/�x�����Uy>��sF�}Ӽ��K�G�|��k�F2�6QiUt�������
����;���zN�@��T*@�VR��?����\H��`���ޙ��,��A��ٰx
��K���76�-���[>-�� 9m�
�-�`�4t�O#��̧1���$F���gv�a��v,�٥N>��ؓZ1�%�a����V[ہT��|���?9=v�ϡ�2�`�ʋ�B�<�Ǖ�/��W������c�>B�"�J[!���Ӥ7l6>Zl����V��y 8A��W�`�}�#J��E�������'`�Y�A:Ke�m�-�w�j�)��^-�lc��/t�(���Ca966�2�JQ��N�5: �x��le"���J�Z��[���PQ[�����i��(��x����>X����v�����$;��?�Ѥ�4gH�F���7�0�}� ��
�D�Y�=
x��[F�W���˄ �V`�/&����!��u�&��=����,|���Ӊiu�Y�nG ����^iP,��po�9J�l.ER C�.sj{�`��:D�;���JD�|����&^!}_����8�N��X�e��F�o]�ѱ!�KѬ�@($-��75�q��"��J��7T�ǧ����OC����`9+Z0'�8-��:����(OU�邉�Sxt-�A�HO��El��+yN���r1��ǴT�����|�J��:6f���
X�צ���`�����Hᥜ훜6j`���܏R1�a��!��+�h��Q�J�_g�������{~C�2�%e�g
����S��D����Zߚx���Vհb!�p#P�V5N���k��ɴ�q���bǼR�%]��kDx�W%�/�����8ɣ�΃*-n[U�ys.~D��X�A��֨^�x}E����1.bZ��&�"�}<�ۡݰ�ztV~[��+�E��~�3�	q�o�@!��h��%���n���q���V�}��$Nh	K�qg��M��
�>L8������@$i �X���!Vz7h]���H�o^�]!R��VPp��b`�q�I�d���=��#��׵>�>��('|��@ܯY���GM�9�QAȃ} T-��j�R�����i0�ڨ�bM����K���!�Ťp9a6��)�Z��:�v,��_���sh�	(�}
m|����-����)�6?*�S

�0�����7�979	l�%����&/�������0X��W���K�<0H����s�z����s��	m/����m<-ι�%�\�B}���m����E�����K�CL��y#�ȥ�����k0.� ��󁂴�M�f �jw��Lx�1k,:�C��HZ�̛�
�ȷ�5�*NSA3�Ed�>��p	R�!H��Y�������ZD0�ٿ,���
���ADk�8O��ULD71�+
���o<3���kYW��o�;L�T���۽,�dE۰7�D��d�Ak�)Z]�V��o޳uĈB�+.��N��<
�uk�N��,ڥ���+r��Kc�K�Cڮ�n���l���Ql@#&B�l]{�a,2�b}H�- | /�,���ZV�T(!8H=�U��,Df�1����lϤ�d�l�����>O�������쬥���0�u9M�z,(�>)�[��C�įÃ�5��iʔ\�u��e����@��EJC�Z�o=9ߺZ��s��*5���w!'�7]m/	��F;\���'�����7��i�O.����0�	S'P���*AK��]G��縝�B�%��:e�so�$���8z��@��\
eN�y����ѵ�	 D�h��Qz�w��9����)	��}re.�K��'%�p�%n���`������w���S�&�6ڇ)y��J��ic��;���|�l��ظD�!�6��z��R�)�����P$�nn��h�d/p��>��3͌������D�]B%��!�W��H$�,|'W�CR��_��#.��?߇�\���AH����?�����#��6)Lg%
���h٪/ן��ӻ �1$=��No���+8��.=
B��(Gx�s���Uc����pʺ��� �]��KK�4l�]i�m����t~R���C��O�堛�o�x+�w�J�h�l[�׈12���\D-����H�p;u�p�K:m��-��"�Pc��\"�RM��p�.���@Q@8[�F'�[��+TT�6y�iA���mx�'��n~������v�a�8��j�_䋤[���/�b82͈t���V ��,, �A@P�ͽ(�N:��6
U����~P�x�)�t�e���b<q�*/�}�P`�S�p�{�;�1��kph�����g��@ё�5�Gw�����h�kQ?��@Y�z�_��f6MX+�4H���Z�U<�$�?b�I3OB$
��A&q*�1/�n)�JU�g\~�=ߟ��K
��������&���.ⓛ�����Y�(�����=��=ue����Zɠ�cGa5�9S�(%q^A�'�}Z#�U>�kK٫�e�}�˪9O���e�`-��T\���&1�J��[������Lj�TkF�ߊ��`J%C�X<�����,[%���>{��ա �z߆�l0�p��xh��Y��ܭ"%���A'"�S��Dj�'�P	D\��� fiG��9�����G�kH��(�����S�OF(�J{�x!�H��Ӗ�&���\!v��'/@\]x�Kp���~�t!ۇq�/�y��n�R���W7):��	���j{��#~�C+��L�4�
q.���4\=��� (�ō<�lc�B�+�8w���O�Zr��N��g�
���=�)��G��s�]g�,3�*��d>]G=��0iAŧ��r<��?1�3`!����-Vm��i��\��F7.��ѻ�,���7Z�H�hjz#FD�iN��^z��@�f�1m��K`A�B}L��sާ���4�L�@���n������%
�.�}z�b<��R 
$�=Nn7��U�J{���Ϭ ��aT����^��3�HDX�ג]U4uz�����lΞ�|_1��V�+��D�f��%l�i}�*�j꣟>��)�D�Fݲ����a�mǽ�
O&#�\��z�li�u{HHV�'�(C (i��B�U�]�J�m~�����պԇÄ[��S�T�\|��)e�Y��eqQ�mJ�s�H'��w!
��e��3Bco�qF�7*m�1ٜ��K��u�����Cw�/��hGoYcL99�MpO�ڼ�-5�"-s�����y!V����8;��RߙFݝ^^�N�f�5��q?�W��@+za�?�NtO`	̛�>�Κ���dQo7#\_P�i|�VOB��B#���W��p�[���޻Y돆:�.{�r�Қ�Ɩ^�w��� ���`��	�Ięy��z��u�����
�֨�f����=<6��M0c�,�gd/;�5�2��D��FA�>�lp&~�����y��/��ʧi����˄ ���;��� !�!A��?��r_�܊R��^Օ���+-������N��r��ג�}�(� �O㓃\I��Q�<E�vR;P�[b9�Iav|#������y�ݗg������� ������f8��F����Hd}��I�(�!܏ �d�C�_;���6'��ұ{;�f4Q[uu��+��Cl�I�?B����r4��e�0nߌ`k���P�U���%���P��8�)%��ZUjmK�Bo2���q��O4IL���pUP�mt	J��kRm�N�&@//�͏���7���쩝jsXm���n���ci���Ag�Æ�W��s�r������6�z�e�Ƕ"�-��Y���d��g�+�>-��gP�v�<'5p,�7�.�)�*-�/0`��T��I�$��3�|*Ө�)J�HE����Bk���q�}� zُ+L�-j��['&���Bb��@���CwM��ÿ��&ʷ��a�V��9?�;�QfV˽W´�[D�H��a`��Ml����1����u�ŨޜV�d�&��Ty�1�b��=���@��I4�p�D�)�������z�����a�%�4E�G.x���DE���Ѐ�0������x��Z��=y�9��
�ߩf
�wNϱ*�2����q�@�Q�8��3t�
臓6H��?��-��ҋ���N8��p��]�tp�W{M��?'k�<��'��p{8pн�bnˣ�>*��}! B$�/A�a�?��)�n<�2%�y�Vqɷ���y���v���ڐ��N�������ݒ/o���7������K�-´�!?�ø!�ä�s�n���1Y#a��n.Ό��3�d��T%fF;�t��#X����+�y�f�Z���5�Cm�u㞘�4�u�Q�Oz䧣��?�{�N&��kA7�a����^L$�[?8;��Np8>*�Z�@�+��y7�T��ȿ6�gq��WU�w{�܃�.��j����P|z�W�8�. p�85:����P�÷�,�s܎��V0R�� ����G�%w}ޢ�W|�1����;Q{l�Ա�CM9�ߩ��iAw���"޼��3��j���_ 4�צ��zD^_/YQ�h\AgܫH�`X�	�I4%��.�[�qܗw��W�9��cT�(���mG���,�s@��~7�Q�#`�\������~x���կX_#��d�y��^��E��H���d�4����E^�G{�X�����A0��O��ke�Ʌ��B��m��(/,!�9fG7�AwFR hQo�8)j:��(��{geB�Q��n���T[��Z�2 �}��+�	%�VOΐ̈����4�-���Y�6bKP�ErØ� sa@9[cg�wh���B/���KK�ɕI�"w�&�ڧ{�f[��o ���"R[7�K7�!96`
&��u��4$2����*x���כ8_r� 9'm_2�}0�>��5j�$2��y��i��F��K#-L= ��@ƮV�V�8\P�:_��{�z��.v'嗄�0i.�=��eo�wxL���+j&��='5g��<��(�2���������uH�$���\�/|��<۹>�\��:^�F�u�l2��|��-��4��:eIS��w!P������y$�3���އ��I��s��h]׈L&��d���7$J�gʓ�qǶ,]eQM 9U>a�%�5�/��iɎS��p�1�n<A�$������2;}���+�^��_���U��[3���ii
m5
y�W�U�_.��,�9A{ΏCVC�ER��)O6x���$PD8BB�s#�E�J��Yg�t��9&JCK��uQ���~5L8~#�a�=< ��ѓO��UN?�H�t���V�<4B��	of�5���qP����k�hnT���V�%j(<�����K�
o͓��	�l�qZV�a(7B��(wo����yw>�*E�xf��(#W���}�\9��V��	��'��J����*_H���������&Ud�N�g��>���O�8����#�@;P۪��}�s�~��ޏĥ�6P�\Ed�p�EA�j`��cpvD������.5�Q�3wM��Y��\Y��XG�IN���-M���B@��z8��}p�^X50��Bg4e:_�y
��P������$/�e��5�'�h�vs}�tc��i����[�����7���fx8�K�X���ۡ������P��
�؀��R夕҇롂�'��U�����q�2���/(�XW�X�h�Z"x��o��;����=I�>-�v2�YO��ͻS��y3��pjϰV6����x��Yd�'�J�e��\�5A���R�+����F��sre�]�� �Ǣ���D���-�X�|� '�/�pJ)v� "�n�j]��$d��AT~���$6�=	��h�� v	�Y��Z�&9B�F�6��P.�X��t�JdP3y�%ו��&�S/6�P��i�*ztH�~T{Q:�?�h|f�[�����r�v�V����*�OѴ!�YN�M�^ɾ��v�L2�������V�2���'g�A{����@g��~3t��(�߿���sY���w��=�"v5��͐7��V�v�N}�߱�o���Ŀ��Ӥ:@���"��V5{7��K���B��kS�$t, �HO�1�(chL���6V�t����s_�25��E!��7�b�uVEӊvR��
�$��TW�Mq�[��Ӥ���jk�����9YB(ڜ ���2���{����s����=��⻖���]MJD�?"���Q�
%&G-L��O�?o�7Aq�jܛ#	�U�AE[�䑄8�P��?�'�@�n�^�7�'�j��+fN��0�VЇ�+O�/#L�o]&?�y�T�S�￈'q�U�'�����l��ԩS�VB �`����w%2O����Z��Q�F�:k��@;�V6��*c4��ْ0�E={#�4�~<ĸ�H��ٕ�e��P$$Psߢ�\(7�Q�S��kqI/v�fڬ*��%ŧ�LxG�[��Ş+�Wt� =vl�Է�?�!rs�	,bj�c4�J���],l��C[�l�fؖ��g,�-�]��~c�&��)jp���+5�v�<��3M��J|��]��lM��o�?yK���'�@*�Ҷ����еG��9mWF�h���>��{�T�8�Q)#)�4u�K7<;�G������kl�*��ی\9���c��W�cH`6lܔD�`���Ō�&��Y�� �V5���=��"y:��B0�ý��Q9��;ԃ� ���IԶh/A�J�mC�������UI�S�7�w4g��)u8��>�n��1���Z(-�(�P}���p��Y���	��_]��o��,�����@k@��5W�B���>��P�o�63�+q����W� �;r�S����T�7�[k��h�D�&�H����IqD�!5��຅t���:Xe�����LM�v���#k�Z����V�����
�+lJڧ2i7�n�a�@�WW�"$���T��F]�|����$X�
���i9'qc&����5���ś@ޢ��fr��C+d���?nd�$Xڙ����cc,~j�ii�Z��Eo��P�pe%��<)�i���$��eJ}r����20Ⱦݸ���^���p��c��v):�\��?���߬�BA���Ks��Z��s�y�Sir�~�̖|G��U����]�-c�� ư����\��1�eo�����*�.��kJrBkJ�#�R�%�eƯ��i�T�GC�UU��V+��DG���ӿEQ�[��}�Y�)ȌG�z��0w]�m
aN�Ȗ�Bȣ��{��ژ�@n� Y����T��o�E�TG����-z�.E�8���x� 9(�,lY�K�,�)p�	TCp�M
�a]���tJ�_��k��Ww�D[MÂ�f�51:]��Xn⚴WJ�;6���Pȳc�2k�[�k��)�Mcp��yp�����2�����Bd�E^���&���uo)5W��c�K�����-�Ϙ�rn�q�w�ս|r�sB0D��|�6Ed�j��/_���y����ƣv��ұS0�*%�=��Hw���B���Ҏ$�.���,�	�}�e<AQb���ā����_0+�!Ǽ�:I��>Q�F٥?AO�FS:떈+'.^����I�0��| {(^Xy���Q� ���<Z���;9�;x4���Hh�f�ўBh=�X��� �p)��l4'p@�e9`�'�}�̀�ą,t�66�;���4�vz^�tW�ԅ�:!Q�����J�8�ς���mg�N|�_1�~6~X��-O���K"A#ur�fu���ns�2�@�$��
�K�Q�fp;��KS��I$��"ҝW˼wJ� f�:^Nw�tr�Dڿ�jAr��өe���c�H
H[xB���"�ҁ�}I9��B�<?�#y�ڶgMb�`��Qs(��S���J��˵8nʰ�2\���훈�@��fԏ�=AG6�q͝S��or+��O�������Р��?}'�I�c/�N�� ����7$�uwrq�}I1}��Z5ѢC��,9���Ԍ{>z��,(������k>'MC[	�s7r�Jr�=�St$XxJU��tQ�D*��4߁��|jq�����Қ/�F2<�04}�o�x�^��
լ��;3	bd&��L���*��8k$��2�M��JsKrz_w����t}. �o_[f�@l҂�C�Pf��+*y��6G� �{u�,J7�R9�1҅=��&©��Q�I�l��fzF�$�j�[Y�8~d���~�]�u�1Oh���q�	l�~mu��g��5̣��W�&�N�X�d<�tݿs&��(�F,+�ϴ.�8��l������@��#kB�2c^�e/$J�y�;cHM�� ��(��b ˧�E&�p,�b �q���n�>^�T����I1��ξ��)Ƽ֓ip��gw3 ���^yk>��*�q�7��E~|� !���T^��0���B�7w~�]sD� ��n���'���J�1iN��,S�8�R�oc{��(4�l'(Hv?�A蝨1���Ռc)��{vp	�}�3~�ϡ�[-I��6�}ڿ��K��a�!���c����#�y�}��}_{nڇB`� �6ο����<�R�V׾�`p8�Uy��c���%U"T̕�!i�Ps���[�7Y�ѭ�2=����������~ 'ϻQ|�O���"��?˧Zi5 �ܧB�r�C?�+h���{���ڹۗ<c^�
�4�1͝�z�D*�?�?�#�:F� h���r>o(��+:E�H�F��'�O��?G�4���37�6�hzcP�<z��eu�&n��[�}�:( ���$_��^��a����S�A�������f'���b!�ߔw�"<�>�s���2�?���`L�4�"A���K���
�"���bD�¦�ݚBz�1��?L��ڊe�5hK0,,�'���1x���p�|s�Z��FG9�ҵ �L�f1#�et|�_�WTƶ�-�2�FСM�6Ŏ"d ����;jɈ\��>����d����l��,u]�ѩa�0�:s
|H�a�'9��\fG�#]�V'��hH7᩻ѥV�z��DRh�-���^v�����I	���n 4�E������+�]�����-���L�o.�}
���4)p��J��<�i�&%��|��k܉RF�c����/��ď����P���YC@q5>�$��u#���Ve��]J���i��J��Ұ�(�Z������K:K���P��M�f��#.�Ν練F��8VD*�M٘1����mQo{���.���� ���k3{D'� ��4[�B]AC�q�.7@���v�#/-h��tW�����-�� �>�t�۫L�x������/yZ��ܑ�Y�0A�Z�O��ݐDxIF�јK�:p')oU�z�PX��U��Ij�񁐪ۥ�]x<.Դ���u�(Ք�b�8|DB
�d��3���ʽNd��%f�_̑J�;�q���h�N51 }t���B0��������u;s�5�E�&�EfP�k�F�N6�J��}KZ�g�P���nVx�T��khU��Q�V��(b�C�k�7e�t�=p�,��,�<�b~`�R�e�
��j��\Y�+3��=�SL�C������$imq��PAn�@�Ѥo�?�&�A��m�X����A�i����ϥ�m_O��E�;B�I|?��C!.�%���KZ�0-�� �"��E�_�t�Q>/j�Pl���:�^��$f{�%�4w����d҂�~������)��P�釤"�%�zP�o�x8��F?�A\�(�PH�0A�m�1���ɝ�~[ea�F%j%�h1��H�G����~"��eư�pXKF�R|ɳ��H/�=� VK){���g��Ro�$K�j�.��2de�߮��utȗm� \^S8�Ե�2�˥����N1�n��\��R��pI�q�¸��$D�X%ޠ39=O��7�M7�mL�,����s��� ��[�{��G�d �o^,?�Sz�_Չ��2AJ���R�Yǟ�fms��;@���X[�H��_<��Rd5h�nXN5tP܍�eГb=8dh$�޹���R?dt^T|M�h_����+��V����-�"C�Ƃ�W�����Bg���l�������$����2{�4�Z��)��5�`�b�I�}�����[��qX�M��ŉ�f�<�oɎ��ݚ2=���ns@�4�:� f}l���1}[=3gk�U�Ơu�3#"��?'Ű+]@E�rd���D�������1�-�6Muz���8�HTr�(: �cIP<�W�Ā>:���"��d�Ov��f����~r) �S��dD����-��$��2�X�&F9��E��/C�F�y�(#�qؖI��+|���,�-��į˹a�&��W��.+nv�Q�qΡ�)!�׋���{C;��Ҽ^3� tJ�u�D���&ƚy��p>�1Ln���l;���'N�%4T�U(������Vt�\��e��֐��E�9�@O#�t�#�e�Զa`iO�g�-����l	0�G��?$'.r�f�KK��˕]D��/4� ~I#BM+aP����C�w�O,�����Y�����=N��f�8���+���J�C�/Oj�c�����5-�������5y�(���+P���j&�dB����
��A��X_z��5�'���,�u�6)&��,SF�����w��F����]}#��9���Ţq7U�P��q��^�!ʬ/��)�&-�Z�}��7٨��_*������|4��Xg-0�/(��M��V-�k�v.*�Ѝ�|���Z8�G��{B��Q^��̛7�+1n�4���k���K`|��
�3�G8�L��E|ugc0Й
��D����}�K�`���\�����]��_<�Сy�$S��0�a�q�&ם++�/�g�ɺ�2L��`��ԕ��8��bƟʈ"���,H�@�1��3+V���;<�e_tw�+����B��@/�V���%V"�Y�0�V~�ф�[��cB���O�F�	Jڟ��4��O�z�sk �#^���߇`��08��b�C��ƶ����UJ�亂-�Ď ��#���5�tr�R������O{������!�򕾱vI�N��y�+�xa���J9q=�'�X>&�Ew��s W��V�_Jb�W��~�2���"�FD�>�*�-.!�{f:;ē~������r�4��b;lS$q�O�͍��ݽ�M:��z~������*�� R:������7{p�?v7��[�z��u$�`F�c��Iax`ܢ�t^㴇Ǆ� ��n�8�0��a�1Ն��.�m�k; �M��ma���t���ƪ�ߋ�.��);����3(s�㜝Ⱨ�kg����3�Fj�~�$��JT��	J��Yp+n�Q�;z���	��Mӥ�Yв�u�"�3�-β�m�%0lH�ߡhr� �Un3L�x<�,-a�1 ��nA�I�P����q-@)��18uF[��$2�7Κ�+�ׇj�,�)3�<�B-h���4ǰj�/����_���JI�w}�>W(<
���&�0y��:���m
�Uio�����$Ĥ$��
�~E",��Z�>{--�-:����@Btn�g�]"h���;�h�f���U�m��;S�(B5�h|�ۍ!��b�W)�� F�X�c����\�Cޱcd:�ldKa+xe6Ű�X��b��N��wtrό]L1k��S�ݝ��E}b?�A5�a�K?u�X3@�R�Rk��)�Ÿ�'�L\�z쿝��;�Ȝ��R�d9
�:��P5��5F����WA?΍b@J��+�SA�zU*>
��1�4�|��إ�'�lX 3x/S85,T����(+�ɫxb���-[�ً��?�M��Z��u�ѳʰB���)�xu$�ش��GTa�������:�K`�=��(�$��!!w�
ݯL޷:�h����J6����H���)�ߞ>�����:y! ���������Ɂ��U�"E¸n���ȼ�#�Cp�)m�a$Y"{��/h/'�H��o�B�R��b1*��O{*,L�aK��of��G0��P+����O9�i��z�U��c��+?���9��@aQ�M&xg��v��Y��G�ٵ:������ї��+[Q*W�X�Q)� �\�����q�px���I%
蕩�RF���OZ^����ff{������C��;@I�tXL=mLߕz��Z�f�9bH��/0} �Iy�z~��I"��D;�FCOݶ�l�3��-�h��~j�hr
�/*�г,���<����G+��c��Q�]�I�S�M1MyWC<���72���$�6%�d��'t��ǯX�'�vO$[T���Q���L����`�}��w�z�춋k)�J#�~	D�}����6���I_��ڍZ���T��vϡ�-��>+����:��b�?[E�%�Ha$�Z26�xQ�>�_��g�����C��D�}��p�VcXU,�3���5����^�8�j�G��c�%7D��P��/�$_f9tȮֽH閠
�������������n�v��#DT ��F�}dN���}�ӳ�����#XZ����(X��MY�o�5A�HH)y���S�Z�ڦB�#��=[Q��e5-Ux���H@�١������1L�J�`��E�k�"�S~�k`�b�2�/ؐ��M�����>� l}D��F��M��%�LR�*>�؇�(I�������Ք��6���D���$��[Cd!�i�w�1��ӟ72���ƾ���ۺ��Jδ���xk��������\Q�&�F�1�/c��6� 5wk|����ҐS��3EE>������d�P�."�G���������a�!oc�/:'i��O( <MP���]c��:�#����v���u��j�}�TT^�5U�v�ׄ�'��֚�����#驡X;QT`�峧\�Cw������'}�)�P�9�W��ˑ�m�KG�2�q�����*ۈ���X���'��N�����a��N9��c狪H�sp���}!�j��-mbF��7�';����܅bC�ȭ!aɫZ0�c֩��xE!V�yCs;}���١�^Gl��՝v���9��q�O$ѽd�&�:F�&�Y<��@�H�\�r�3�*��"�
\��fK�z�S�z�|�9���?H�8����C!�ۥ�0
��i"���٤���7�̺���f��5��©�,��6f��qY焂�c�TeK�����~�P_��f�����]ҏ�b�o�g��_jQ�=�k��4����ZVۙm�ˡG4k���T+� ۨ9eC>8R�)����,�y��o�Ė�q��٨g
V�qW�ÓBr #ل0��KL��b��i܃^��M���ܱ��YO?0�+{�
�%�
D1�ն/v���B�A�B��_��CB�f
L�'֕X\ky����u41ه��j��t�{����,��ݞ8*h'��*YիwcN�s�����5�Cv�~&������wʌ:z�#~�ch8�W��],p��8��R^�gX�jKfW�7��"Q{���:�����X�1���-3�%�*�W�Mj�Dg������tׁ:��^��6���kA*d�k�����A���7G��)%�އQquǟtx�������G6��t�ܙ�Y[qF�B6�>������}��uF0jyLMPq�wv�ԫ>ϲ[-j�e�6�%�4�Bj�a�f�������,��Aw�'%Kq�?�p��J$%p�ء��T����=$���p,���!6|�Ԯ�]u���5�]���7p
��L\j���vK�S<KZkN�f`�4�Uy�r���q�=}��=@��'>�7�0À��������33���;��9��Ʈ�cx�6�]Ճܫ�*)[�6'^)��< ©+����nfl8갦�ٷ�����O�ƈ�Y��F4�����۳%���g^M�@��3���_ԙY� ���n��H���d�����w��n63��%^�c��_�~S�J�Yx�Z<V��ryF� �9A�L�%0F�O�^��d�$"�>���ºd���4�ưd�xv��p$k��v�P�ĬLѵt>�&� �t���J|~�����~������W���omE��1�h��e�GP����P�8�3P��6�
���Q�=M��A�$�NK��|�k�5�'{��8o�ˑ��O���$}tl���	ש�٫�_K1�R�����\4�@.�#��pm��I��	�P#OJFTM�S{O�.#[�n	�
�q�#說��{�@����5)��^K6�MӮJ�N���gJ��w�����ٰ�������T-�D�E�@ĸ>n!E&[���0�V��RF��nT�{ci累y햱%S�l"�,w���f:]�

�a�@�������l�N�<;#�k�.i:�Wg���]'˴!S���*d���=F��7
���y"$0���&AN	=r@6���ke5����D����݈�_�K�f�{Q�SHK=wp�1)\a��11�W���6�k��}Lcp]H�7���%_����̞.f��^½��
�A5¯ �J�ڟ<>`���XZ�/��U�6�d�ATݘ��Z�C�pM�4���NU)!Yƻj[c8xU�1g�0�b��s�ȋ�q��+�^&��: ��	�M ��y��y�����q6��:g\u�db&�+���	�Z%�3E�M��{ƹ����U$V�7�o�n�rt�	�]�ZK̙0^�ďpl
C�0�	��B��S���[�]���B�������Z	����-�
�A�U�T��]�~�y{��S��*v�X/�~i�;_ك�=z� 2�n�Q	��"�[���%zuZ��B*ڋ���&9�uET`����:a��6�x�^�Vb�ӵ5bVS�W]A�|Bg� ��|��#�B ʥ�*j��
P���o� L���?06�||���f�y�Us&M�s����m�/D�'���U�q�8b��}/^`�>xR�	V�v!5��3A�ADg�D"��p��j&�?�>z��1�=��\�w�KG�73��Mp�E	���Y��d	��e�]�ۀ�a��<��H�M�k�%ؐ�t��_�����l|��Rq{��kz��G��wh1��}E:���fQ�@�G���
��c~sF���!e8U����&VnYT.��,@��`O�R��M@�N;�W���i�F�/�UEP��{�;Ϻ�����/9.o�M��s����]�"⭒��ڦ.����Al��U�U'��_��|[�H[�A��H�m�B2��Ӂ�B�@V_�j'͸h��!�_9\�s#c|���!�u엘Ú&�ɞ?���;����d!��)@�8���������������:����F�4�1=k[@}��P���_k����ŇqQi� CRFG�	��w��~��	��>���F�a��J�	�<[�ɽޏ�$ڒ���=VS�����Ū�i�Ɇ��=�®H�����J��&^20���cE�Ϋ��PR(j�	!���=A�p�j澑��=��L�`�[c V֦c�������μ�ep8E������H�O�T�٭x�p��BqX�d ;ȝij�>���wG���6:a*�ʱEg��X��3�{�M"�j�J�����I3�5e�l�����7�B��v� |��*�M�*Q@t��޷Xei�V_�C���;M����ڑ_���0���BF�Y�&�ʍ�ߣ;,>�Z����oy�B̀�:̈F�`F=�R�����s�'m��_<���e.NJ�K�;� Ξ��8O���떌}t�~X��b(�fS�MIV��
7S/uT(�^y/�Y9�B8Xߕ픑����M"X�d�4!UpQ>p��m�SWw� ��K�Sⷄ4Ko>Gy[���syN�'�m�-e6R�e�:P�&w5m^&{�V��v���@B�u��r!Էr�ToE�p� ;�.OT��Y̔Բ�1�W�ϓ�4�kǂ��ʅ �2�^�:=����f�.�+�'i������BM�}��iw��ʭ�!�`��}�:8�X��x�+�+Z)y���"n��~���[�z����F����Pа��q2�-�
9`�V��5��d��W��>}7O\u���朐蟍`�'*�*�0�x�?'L�z�(�kX±����X�V�)œ���%���o$�Dd����
zVЪ��`�j��'kP�mI�����0�i�L.����[�#JZ�ju��Yu=�;�7I7�Y�(�"v�)g览�����a#%4��i;��g�pJ��H�f#�,[��1�y�p�n�"���xx1e��I߿o�M�����)�������J�-!�2)W��M�^7qw�:�C��_���ĥ�fR.��A!W�9� 
�3i�k7N�]��4t4�nD!�+ݍ�-^^�*�(䦼�>�`ji��v?a<c5�� 2�&�vc623+�j����8�Z�@�]p\�I��@)V"�����R�'Ҕ�M���㧗�B'}�e2�=֩�c�jo�A/� ؐ�&N��Iy�RU����.����`�X�iYx�����f�'H����jdP+3y���\��`ǌ�{CLp6�N}gB� ��K�c(j=�|k�}�GD���3RB[�7��w{�BW�nd�ˮ89���6(w1���m��1~���$1¤�{����u4�f�3W���%2r�	��4��c"��>����a�`���ҳn���fO|.�&�{$2H���.k���=?:��� ��#3e�	lrŲ$_�	9�L}����y�tQ*�t�^����;��)��m���HN�N�X��+�tO�cJSp ����>�����{s�v�����3�MȞb�(�K+�Qtg�z�#��~�7�+K�����M^�Ų
��ɩuEB��R鶇r.���bI��m1����2�T�ɩ�ʘ3����rϯ���J�螤��?M�����>Mwð��{'�,���!�- �*}�"K�'�B�J.�Ӏ�?��AB]�7p��.[�����&���x�G�cZ��/zy(ퟕ8�p&�k�=aR<A�x��1	�v�H���S�c�F~�4�3����UW�J"�E�KԦ�UB�!9{��?�4G�@��k�ɰ����%}���+ˡ���m��B>��:����� ���`����Q��������=�=g.~��t�C�Ƥ��k�Z�n�����=:�_1x�ds�c��39�IqG���S�}��4�s]*��������m�u*X�Qf��H���z��8�:HZ|>8:���"�H%F�ΛE���n������`�8�$�CxO�"���{��@���=��ۧ瀴���S�N�t����$�k�,�v��;{��T�t��s���n(�$��I�}П��p2I2��Sv?S�)~U>��V��g��!I{��(��tNb'WC�T���o�j
��=X�$w����qU��ɬ���2��0��˛�O񪢉Ԩ����]�90�-X�bN�	��G��l�n=:���RZ��ɻ�:�Ŝ��(���J�9o��br��;f!�G+�Eo���qb����uԠ��}|x��k�ȝ���g���ym&�Y̫ 4u+BpP�8<qR�ŋ�(��FG���!?�t�}�pϟs躩�;�O,���/v�����/�l��ZeJ���՗�v_���'�O
e��C��T��� ԺK��0� ��@s�:P�Tu�|sL���X�i��#��uf�
�
*?A�)jV����1{�;�  S��x��);W~sӻ�{�3{��bW	I�Ŋ���u'�����_���'m�~�\�ǐ��������<�vYC�{��$���Ddؼ��}0�D��������'L�'Ҳ�g�Ƞpi�}1)�St#F�?t!�84g��B� 4�F9m���#)Ҡ��+T��[�8������MҮ�����^D�8��Y�6? a睲H6ь\�9�z3�T��t��K�C���Y�U\�~\҉�j櫮LR����t�� n�g�9rUt���CӧB����,	���52�!˔�.:�,��$�?������&y�%�!8�e�B�d6���`�*Hn�]�ک.,��O�9#��ղ�7�������G�^�az{��0q^l��= �KQ��T�\�����ؙ�@�R��]�tY��b���!b�W����Uɕ"1Qu%+?��?�	fZ�K,#�44�m %m0NL�kJ����BH��q�>34�Ɖ{�"�RO��80d��W��Q�c<TS[(o��G�;�_{�wOki��W�����{��桰[l��3lg&�c���g��G�8��3?�����~�<c��,�4�_N�އn[w�	�3'�%�5��o.;	���f�%��)�?L7LÌ�MǙg�݇'Vޣc�S��wԊ+���?�M
O�t{�����l�>�
q���<H"��rll����5$j��AE%;~0��u�6�����A�����U$r9Q����W'��7�����A��2#%q6����@����*�D������I>@�M9�C`	6�3�䐢Oϝ#�#��k�ѣ!CQ�)�Q��!R�>���Mc���1�t�ǳz���B>]��~��Ѳ��_%K�"�	"<��y�K��t��0Z�[}����\ֈ-3-8yx�&>��'�"(j��Ko��lK6��r�%��� �XcB��F�,L�$.���6��8E:Tv/)�Md���:�%`��]5�.n�@./�f�v�)�$$kcS{�V��
��3���Or�6���_�]��u�i]#�X���zL\�.���Hy����W�y �G}y,^<��s
L�X�>�%��A�W��J�6��ɿeB�-��p�Xb�\�u�+�<&ͧ�J��Z�ɸ���tB+��[�1���?���2�┵czG�	)�ۛY��\CL|��a@X<���%�K�}�u��e�!ː�/�&����P�Ąޥ2��d��� �pŖ�2R���3l{%� j�p���=�0��=��:8�uT��o5}�@�p�C+��/����WH~� �Q{l�N[��L�01���z�9�rkԭx��޸�!0=��;t����Q&m��1H���P��e˚yy�q�
��9�C&�xB�,��>0����+���n�3�mj�-+y�������r�g:N�`�����bto{y���������s��QwgM�$@vX%�5|���ye^j�����e3�o�R�c��s_��.YL��4kp�����D,��+2(�ƈ��rꑓ#7b�ri�t谚����K�-հ��YE]r�꙯��,e?�����&��27�����x�_|��Ąo��|���=]���m�6׫q�d�I���e8�D&�6^ mL���ݽ,�&�Y+1��C��g����|�a�d2��a�����S���I��5�����}H6���Z+1�S�$�{��23�8�n#��h�0�b��kWݱ�rO�k)8h��*/˫��a*��_Ez�?b�1:wau�EM�n���Z
��Ʌف=��u�D����	-\_��n��$N5�tlz��6��"��<�$?�IO/����Q"��5sss -��U�R�ob���x�޶���'N��oD1��p�ٖ�@�܉2����Z�Wp��(\d�	��&L���<��H�TAm��@	}�o�Y����(1u�����	��t�0/�|�� .���,���!�8�ʾ��LN�9�I�/�fՔ�[%K�/�p3�Ƴ{���s�9/M�I<�c��_��/q�ƛ���;�Ö�#���JTnNWԂ�.���ݦ��TS!��������i�4��ul�e��#k�˴uC��tD��R3�K񣻁*���J�������dp�?��\�ҭ�i"��s����w N@f�z�]z�-s䨭��e�e>�}�4:�9&���3}�σD�b]*�O���iǓ�]N��i�0i��kQ��~9�jg%���re�f(�M��v�w�SF�
��6nܸ���ɏ%KDof��"�?��U���J+���K���#U�
�:}`�	-	T(!�(�{E�A�	M�:�3W]}Ҟ�)��f��\+?V����c/z��W"�LB���Esa�M��A��Z�a�xVZ.��ݣ}3��/vP�S%[y&9����.��m��(tAۓ��f�Cү]PZ��D�yzP��C�ZM��Ko�f5��ґ5 �Z�s��Z<;"q+ݼ��*�f2Rf[d����wo�ū;]�E�i1W����v�(�L.w��OBU۴�N��rT��{�#��j���_ǈ�|�q�?!O����J� ]`�J�mvؠ�2�J���V���a����Ԛ����u
�(��HQ�g�s
ܱ��1���	~@nh;����A_��v�x�[`p���w7�w�(������}(?0kn���o��{��ke���fgp<ݜ�Y��w����B�ep���@v]�3_r@���A�]��ݝ�?l�.����S)�m5r�A���8����$A{��h {S5J�V��X9�Sd�ٿۣ��C Z��Gzv�|'K낔"b�Lp�^ئ���}QWj�%PR3��FP��YG��N������b���2��k��z����c��g9T+���#+��	W��4����/��V:�U)��_�g\-�c�6Ofg?��i}��?�X;Eh� k��<�aO$A�e��J^ig+��0Դ-8Z�\����T�J��E
%�Ơ���V��uI�t��wV-|n^�K�{�(n��k�4�{�A��z41��=|�a�F���P�����	����H),��B7��-a=]tnd /��X�E7��`ƴ+0�5�����Q�+�3%�ӹe��$�+��D�g���0�x�k�W�]//ž������в-���lH�[�v���u�v��D:qo~g��4��,��.̕i���ը��lz����l�Gs�є$d�W�P�h�#̼Y��i˛+��$�$�펬E�e��v�_�@Y!��y�\��ܷϡ�f�)��ª�\_���9�j��|�(.�bl�L��f�o����̒�_��Dh��~���Р�9�ʶ[�� $�BQ�8�'�˽�V���D�ɂ�s,_ݸ;�C@�(zX��_��] ���	 ��ʗ��y=Z���VR��B�F7�~������:��;^�索����0�̎׶J�'�쫾������p�K�K��]/]޲(`W9�M�[��e��������RF���Ě�YhR�8{gIR$�%&�h�q;�P��'G�r^f�;͹y����h���;��u��n�r� �D���r�u���'z�H��^a��C�/Y2�HR���O6^���5�I?�]�[.�=���+�Oe������HXd������|������`Q��r��0Z1G�r�(�����]�cIh4���=Z���2ټ�p�vMs���t�V��� �X(�o���eZ��._h�ȱN�.���e���M�V�~�����P�l��?��F�X]_%-��'�����@i$�
��g�P�yZ��#l 񺩋5�d<R�d�����|mr���_�(��	~�l��Q܅�&	�����3���7�d����vD2�HK��3S�a���־������K�������P��\X�X-`4. .��p�X�{�:�H1����5���S���Rʃ���l��8e�
_'�h�N�:=��$(��:�$f
]кg>�CYCO��Q?:��?$� x!C!��q0���e���%��[��f�<)�x��$E�O%�����0�fՍ�n�:Q��׆�EH��(p�M�������=�\F��g��N�n��iI�%*��Q��9Q_��P'�+5T:��B׶���i?03��3�.B�����c���}F���*ZZ�#`ぃ��f<ŭM��b�%�����s�Ji2b�ԗB��D$%�2�����:MP`!CXw&�$��n��` ��_ý��7������ۖ��o�MPA��_��e.	���j������*�������=LE�o�n�%��}�8:_*f���]'�o�gww�/V8�u��4�.�%.V�z�� [\k���.�.��9f\�[���4D�z�ѷ5���O�R�ے��9p]dM_�~�PvAx9�5��\k��8�T®	�����SǗ�i�*�3ՔM?�A�x
T�Sq�n�R�䬔�LuZF��Q��h��+���s��Ϩ���FV{_	ꇱ�Jw���y���v�Y�*���ɞ�PUT�- �����������S7>cn��_�=5�]��G���r2�NC^� P�K3f���I~:��F��ű���^yd�dPu����U�?�O����X�+&A#|/�5�l5�+��%u��sS��)�dE�v�)�+�Ȳ��!c�(?6�o
��FS&��-����Af2^�c諙��w�n9j�۬U$�E&Y��ZSbtp�6�X�\�1Tb8��O ����V8�����_%|\����BQ���0�a��fh ~�]}Y��qYyg�����I�,�/u�d��PĂ�+Z��qC�iF��F����TTE:Ӽ���4�w�%��;V��i�]S �]����-��gJgI�c�3�c��?�p.��E2�H������q������z4��~�k��h��f�o^�!^;��WQw�$��1j�O~�2��N1�=J�q@C#-�o�X�+O�g�py�G_��/o���<��>�ݴS�B-�(��ne�ػ���	����A-�p�*�h�z��Q�
|���z��ˋ�����I<&vN�g�VP��5�0U�fb�m��T0^-����(�\�sG����3OL�/�+v�b~S�a~O���p�⸍+e�l�~��(0	� 0��f��e�'}��y�����y��W��؊Th�>w�bO7,Ѐ�S2%�FR��<��?����$��/����8P���B�rh���pX[8�3L/Oc#�P<o���M���Bo�p�R�`9��l�Oj��E�ʘ.�G�b��Έ��Y�q8A]46Q#�¼3rY:��[��l��TqN��s���֔tV����؏�:�{�����Tf\��X����7�S��|�����++�4�[����Pg�"��<F.�!~ٿ���E��朦�����۫���M��|��[�k��0鴊RIxZ(���ޕD��E��͟Q]���ٽЉ7��ކ�ձs��Q��k6����� �ytX��'b��X$F�U�<ɗX��_�C: �&�*��s�VI�*�YҖ�G�`E�_�6)Y"kK�d��~�A����vY���z7��;�F׃�Al��@/e[��y�F� y4��f��KP�w����v����_�ٛ�R(ٳ���G6�ҒL.�s�]�|�0��/W��G�c� �V��z�y@�����K7��$�3b��nR!�ষ�4�mc�^s��X[M���2��ٛpB��%�b��#aܛ����{h��#�K��jngF-O�Zjť g��i�]QS< �I�|%O`�{��v:-���u�.9grK������o��V*��T�F�Z�좽`c�ޑSl�M����̀���o�ܩI�ֹ����tu�F0L=�M��_*�����ڬ'�9���JLHB�Y�}:�Q�Q��S�#/S�zi�5��k����w4r�vdX�C2Sꁩ�ra�zK[6N��y�ÐV�G�f�	�������|1�bK`S&h��~0���O^9�p�|�a�YR� \nTH؃�u��"R��"(���NN3�+��=Lq��a�CFW)|���}���T)<��L�j�&����S���c_�B=\~���C�m1tg�3"T�U����<��ªq��Mc���/?��Ϋ0TE�����ēj�k�q�h:S�ҡ�J�P�DZ��
O=��l�L7���C���
MCش{���%Ww��� L��}�z��-��輲.(
D^����fr����t�����}��'GA:���M��-��
�L<�6�v���z��C}�豍��]b���g��������3
�%!��'�[����˶�Iom!��T����S���'��^�W���15!m���&�B�/���P��i�����	cBB�o�LM�,e.HK��������( ��q�1�B�@��Vs�@�WL$O*�$��6Կ�x[>���Q�r@J�z�2쮕&���B`=C����R�M��Q�_>.n0��������-��{����F��X�TX�M=>>�Q�^�N��"���4��'n��U#65�*�%2�§�B-
�<p��N6#�cJ�S�=";i1a�o��4��/I��6��3�v~{V�)���)��r�0^!3�ͩ���E�^�ڭ��OY�G}�+���� �����y�?�ׇ�iW��].H1�l�`�<�nȲ��gs��G���ܥ6�m�v�@��.%j)Ms�a��Ȥ&"����n,6�'I��ަ�*�����f4W'����'~	����[3����؀�Z��
5/>j�.80�`�Htw}�t�)�cE�4�:�m����ٹ~͖�9:�@�lG�u�� L,��J���v;�s�q:Aɝ�y M��C�1�>t��1�@�N��Lķ��v�]������JQ&�+*�Lz������^���֭����Ҥ
-i坔`��m�*�V�sq����҉��E��a��B�L��eӥ�-��X!$imi�T�e�i���4x᠉�wj\u���KE�y���ȼu����.�n"&X�W���fX>l�oNu��V(j��\��L�X� �����Kx���q9�	蠦��je1����)O9���"p��G�t�s�jܔ�5��\d�C	}P�+	�P��+f��iݓ�YB�O�)G�oK@3�x����W1�<Z�Ƈ=��X�|J<��}d���Vq	��\���#�J�Ƭ����ؔƁ����!��ٌe,4���r�TO4�&�cP�d��u�ѓSQ"�MF�#��t�cz���JC�g��;'M4<�Y��=�P{u^7�9ܫ�a��MY�`)z��f����,�������n������y=:��#^pЎٽ(`4 qA�9�{���P&&wW~�}���L���	q�A�^[�����T�RDI~��}��*��6:gnԹy��ad[��k۞(.<jH������}T�}�!+�I�����z���)��Z�I���<~{��0��!97^,5_�ڻ�4�#-Gf�a@*�!Ӂ	6�[��Xe�3%��U@���1p�J$�`�Z	�!�Z�uܿa���z_��b���xwF�6/�zoL��L> �e��gC��DJ>.A�Ay����/r��ڷlٲUco-#�Ÿ*��.��:�|��T�s��O�	��L@zz�c�cX�T�J����Ÿ2!>����O�t#~\[�_�
�*;�6ߎ��5n��@�Z�c�����
 ���;�fY��/$�� �Ƚ��Q�|���X�I��]��ŐU���`dy��Nw���{�v���6k��!no��m̹=����y��;�ME���A*o"���w�4Ѳ�>~��!4�y��z`p/�ҹ�Z�����|�&����\sM�F�fBS7L���:��n+��`W;m�eB!�wi+���O)� 0�`M1����;e����E�;��_�R��2Ն]c-6�-X���S�7і��f���6���i�he��R������T��s�r<���"��Q�GZ��R<a�AKF������Yqvj�1w\�a�\��n����B,#p㳕�ŵf��n�L�W����������t���8�츀�������@�5=��W`3������́s|�f`��t _P����w{c�!�Wv2ݜ[��iӔ�TU:t91㠋6a
PI��3���U�^��~z5U�<�����E+]u�k��p0y9r�"��R�Pd�Ȭ]~#iOV��>���<�a��l�
�+a��Í0kk�|��Ń�h��"W1e�2�fOVl�V�
��t��^0j��t�C�B>SfWD��n�'8m�D!!�IG�.��^4��B�9������9�e:l �&4�s=�Sܓ�<-�Ef#:�a`&Ԃ�#����4�4�.Bf\�V�K=�b�٧Lz��W����V�}�94��	s����1��C�Z>s��ʹ���ܘ�;��Z�[��f���ĤW5	���y�P��a-g����_OuE=K4�ð6�������A��6���F6�(iLt��d��0fU;e{� rZWG������#���L�J���!C|?UPl�7rU���o�w$��i>��8v�h�!��}���i��e5�0n���$�Q>O"W���1X?jmĴ�,���u��Ej̯�����҈�R�g�L�<͏�%���z�	+�)�-.Z;}ѵʊ,D����2�o�ކV�t���Bl��"kB������mh@Ϊ��B7.:<T@�f�%��n�gY�	������1�v�A��)' �q����~��F�	��"�.9G��������=%��k��~!�8��q���Pv���YǺ�����o4j� )r�P��mԆ[��Pfb|���,}���v�@�&�݅�W��������Q;�,�F��%P��,D'�3a�\�ט6ԥ��������j���Q��=��!�2BE�J�~��p$����}q;]��SX���A��rYy��@E�t�-Y�c<I�y��/Qϛδcqa�A�����Οa��������8N�.FE���q�^��M8݌$�t���M?��K�S��M�M�@$
��|��h�x���{��'aM��S�I/�*T2Ǣd��~�.��Ҳ�`�^	��&�Ҕ${�#�L/�Mx��5�$K��'<���z�C��lS�{�k�'O�`·�&�U[Ԭ�9�����U��8���5��3�E�R�8�rT{��\?C�����|�2\n~�y����Կ���{��t25򽱈���C~�����\$9&�2��$ߝ� ���{�� ��gTZ>Vh���`ϖ0r�1��`?��K �w�0���
��'n'�.K�T\���AB��R �Q�V���M١�=j��L��
U���!��@sz�$����}C&�ӂ`-�H���_�9ka��R���7󊻢���\�B��2q�]ކ°�3�#k���H����o�5��>�;%z4�G��-[�0F�����f�֠�}?�*��U��"?�_mL��γ�Fwe<�*Mv��w/ܼ
9��-�}B����R�G	�8���Z)�v&�Z%�����fs1* `����$�	]�l^���v�~�vͮ��"�}s�(=[c�S�ޡq��9mq����2�]�8�q%�{k?���t��C7|��S�A�u�̫���J��RV�u�{b�5ˍ�V�e6�g�S}�w/��6�>%9�ޥv�eP���nz\�2����a���=���P�ngeh��lך
�DS��~	p�6׃�*���9K4w��l����
����/�:�nOF��\���K�A��H�z9yhq��c������'���_�������Ka&s
�oUv���:.r��p�M����Z�a-�	n����.Pܯ�m)0DIth�V�\����kd{u����.����V{ō��9e�������PY��8~�qqo
��.��,/iŤ���'����yhs6����d���Jm.H�����rT\�i�����%�xIA}U�{dTN$��ܧQ�&�4�IG. �	�v,>���m�8:Z&d5�����5�Y��c�C�����-/Tt[6�����`�'�D����%o�*Cc���ZVXa��nau`��b@���$9 �����eR|Ծ,!����.�@���4+�r�4B��9h1�pV����-4?b@أ��z���(䌌�w_v���ܜ��:�O��-�e_w�m�(l�RI�\d�����+�8�<O��P4<��[����d^I%�9*�,F1X�e�b��|�ħ�xSn�#���@�(�>���g�ƀ���׍�G���H�(VeW8L!�V�@~IA�A��Po$�<�7k�/�%�W�fl�j!|����&K�Ԡ��-�ķh��tWRb�����ZVΕ��:ZMJ]P�}*V)#�.��s`M9G���v�o�#>/'��#��fcr����r�zH��e=�%_z�n�P`��b:��q�A��$�R���_��~h��&D�oIF�|g�~��"����c�����}����t��������s��k¼o����+"��OyΓ�20���O|W<�+'΅˸�N�%?�g/�C��5���V��`۝1�v�y��j��-/ެ��:I_�eXnQ3������T�¨�5F2_����'�j͙�ȂvM��Aw��1�r\U<JN�m�4&|�S�o�(�И�����&k���]oR�Q�g�=��e͘��o�H��k���}C���o�>�f�D�A�I��
,�N����-�t�r�"����F�E��H�2,�?k.�v݂HZ&%���xS<�j��1����V@��+86G��+��ٵ�+���w�t��E#���5�ڷ�u.����ޗowMv����O�sK/۱J�R�9�j���$p���/��9i�M��7X��u.�B�o��e{#�t�m.�E�?�F�,6�:�"��ߊK�6�t���b�NG]C"����fct�hpBב�*�h�?VX�"��y�j��uH��J�A�ҩ�Y;F3��X]�B�vv��~��v��/�T�ҕ3��~���k�B#�J[�X�
c>��X�g���9�HF�7���h3�Zw)��1ap�p��Q����~��0��3V�W� �p�ahHҋ����|��=N��K��L\
?�HOJ�������H����c��=� ���o>����b�i��z�*��)�K�������c����lwsI_�T�i�-al�Ϳ�1���|�+�9ۙ����d�XL�g�J��09��c��!2�1X���z�/��ܽ�R-�29�1���!zP�Q��W*,o�i
�l������-��L>�#�;�F���c���i)����:�<�f���ږ�+�AM�E��C_�jͷ��ݓ���h���_N+�D��
�~�7V�녊`R���W`�-	R�y��1����o��Q���_��~���g�a=$���3����a��k�EVj�];[�;�4_�"g�W�[����!���./�9��R	,N��ƫ�%��=d�oJ�Y�}�&��Y�h �䕯G�Z�sug�����o�x�-R]U>r�51��6&<�ƹM)4#@�^p�v��`��~`��?]V�l�p�+p��]??���H#�9��DLO���C��d����:�T9�{$��)���T1��F�g��]�F�.l�*�>v5$����iJ���4�l�7��bw���"��6D��U�@�������M�`j*	}��d��>0���q4�H����C@L�~F� u�QO�!86�b��.�x,ՙ������~ŉ��u/,��=D�J�K�Ru3F
֖�S�D6�-J�Ni�7�Pbq�-΋�{le���}c@����(�WK*ZbDI'6�W�n�ɰC�g]����}0�>�j�'c~h9�b�s�d����P�	T�%�S�-X��2������F���1S ��h�"���B�hB�E�TP�Է��}�#W��(�F���PD8zc�Z��EN��\�TĞD�"�v�\ikK1�}�q/�Ֆ�7*xS�Ϸ���?���/Vi���z(�ˁk�6�R,�"��f����4}�f�~�Cc����[4�fk�~'H�N�"`
��d)mY�����n�!�~���2�e�ĳ�e�C���	��a*nQg_�vGC.j���N�\`��gV7�UM(�oF!�*o�^O =.���&�V��&D�5Ĉ�fL]�wq<!vnj�@�	�'/^�kN�ւ�G"�I|�f���j���Z�l�k��ُ������Q�V����L���|�?�;7���Yg2��K^�������T�a)���";�|�m�j��|��GT��5��PE�L�X�BP�*˚�H�Y�stM�=�!�?�~%�i^�)��:��ߓF��3�Ie[�Л�1�E��J'C�����gW��N��sBfq�h�D��\��fE��QRF�fw�v;�@)~d�ܯ7�a,WC}��Cd��b�'ycc'(r��ܕ亼מ6�4��q��{�@�����1��i~ʗS����1�A����>�&S��+�s׈��c	���N[����cL��C��~�z����p��v�In��!��0��1r2=�Ch�H&�p'�j�󠹽GFȵl1�T��5�cvw|�\����O����[dXJ�s���L{#[�-̷����*��x_ᶙ�6����ǡ���6��!�Ԯ0�����8�I�� .J1c�B=z�pI�F�m`�i	�!n�C��To;?�tiM����8[ 2���&�oRp�H&v����X���Xg DT��5��U<�1�WrRI��u`襫'�XL�R$pu� �&<�(>k|@�Q4M�gK�P8QQ�W;�l�AZ^rJ:�3�?x�ٍ�"��.1�5
�����&��.���7\����`�Hr�U�aԿlu���X����{
-�@��3˺�(,��g�Y̃y�&���d�	�����8�!����7kL��̈������5����~����c���U}%[ABoBh�^��Z!��&���v��d��z4��7P�1n7	�S���>e�/Q4�W*G����3B�2<�!����9��D���9�G���Ҳ��H���ӚR���$,�Г������N��.�<
��Av�ǭ���Ŝ_e����8�ʙ_�-�5��9R1�:R�v5*b��h=q�棨�1�nVi�Ϋ{�ɐ�s^N	T�
j�#ց��K+�sRNʦ�9f ���m����-H�$y�6p��gV��D��l����t`,�l�SF�[�tJĸ1�X��g�J��@���`��!�S%Ĵ�����)���u`?�9��͞x�
��N?���Ⱥ�����6x�K{PV���t\i\�C��L(u�ٟ����ܳ�|H���*U��>�O	�5�Bb�T���l�N��q��:�@u�׃�Ƽ��}4���U�UԄ���p?!+'�j;���E�+:! ��M�Pb��i�i��Z�qQO9�����?����@�u.	����C�`�v3}jU�|E i>FT�3;�5N�X����u�ר0x����,�.��-;dr �Ї#�����O O*����>M�0$�4�/����a_�^E�z����X�z���Ey���k4 M�<3��f�F*`N󘆌B�}�nr��!!�f���K��.�A�g��ٛ���q��)����ڐ��9������E�S��?&�Ja
���B�'f�w=�H./��U~R>�G@!�ߘ*���D�6�{f)11�� �ȓ*��������}�E��wW�/��g'�{&��v��G�_��UZ|q��S�!�Q����Z[�p�zW�d[�Yc�J6�8��!pJ���~�뛓T�+�ծzW��z^�fX��ͧ2�/(Z;1Gtk�;ѓ�Q�\�O���z��$�q�迎�Y�:�:E�i^�1�
k���FF]�
��j��c���"[c�'n-uyʵY�%�+��.�ăgج8
��&⠘��`���&�N3�S<���z�W�94IP��?Ԣ2ͲJ7�w���r��g7Ç�Mu�NFD;�hm����p�F�ƚh��H{���i����[;�O��!!���C(�õx�K�\�@$/�l.�4}�ē�|X�C�E�V�%()�F��#�ƶa�vId5��x�͈NE;u���Ɏeq%���T[~�+6o�s����;x'rC�~/�eu&q!6�����|�mt�ƖeÍ@�����I4����>@���3�,^��t�:X&0�R�_�0[�z	腋�V]m�O�&@"��)���yJv=7TO6 �oB�M�"z�z"���.˻D�FQ�ˊ�j#Hv�B7����T�ZU�p��S��_�M֞ 	�bu��s5�YBl�;O=_@S���?�zƉ�*E���}Z�����z94y��M���Ir��2p��F�VRb�ء/��[�v��b�4Y7@��ĹMP�%��U]+!*���&��1�����y}u�|�Y�/�a��1s�$�B+0`F�n��pb����Ѻ��P��,�j������~�.�aAϾ���$`> h����oY"gY�������ٓId4�ɽ�R���P���D5���Z�ܖ��n���1ޛ9O(�l
���A',(m	�x����"y���ܧ�=4'[C(�U�|�D��&��Y:	��RDh�S�'�2�� �鎧$�y�d!_7�:��{eU�l��
�����<�#&-M��T�6`�;^���X�+�W�_�GtdH��]z�^��<e��ʔ1+�(:4�=6+�k�@a���u]��n��.�����ņ���}E��n@������G��❥TI~�0���-���f���y�Z�dx+3�k�-�kO��n�]5�}�?N�	>�xnU��f]H��E�>g�Hӿ�n�\�wb�)�5_�8�8�k�Q�g�JF<Gv�ȱa����E��М5_�f
�i:2Pw��1��rk]�6İ
��:�s�$`�+��_$�jk|u�Eʟ=`q�5�)��N��)�8���~�D����q=6%�r��#�IQ���E2��k��/q[Z�*
Q3>�($:)(�f�L��}X�P݌[�3Hi�[qZ�����,ed��� ;�?6�x��5��{�v�1�i2NB��B�Ac� ���+�9� 7��k_�E.�ח�Pb���.����UARc��8�4<!3��:���\�0%=e���ث��
	�r\��ry��հ��:�f]��6N
mU�;K(��ɂ��t
��a� �G�kx�O��0�uVv�5�Vq��!m�0�y�?�ҙ%ϭ�k�w��ˇ{�<~�E�>;�����t>W���4R��R89�x��B�@�T^���@� H�n�^������4�N̡a���+H�J��Mt[qJ��@k_V�����mx�[d�`v��""�zL���P_�_�Ze�y���<����o�F!�o{p>K�<�Y�th����|)#UH����*�4��ct��[�1���ͪ�B���U���zQڎ��D�ӊ��\��ŞEJ�m�V�Q�hlWS���uL�{	@|z�7B���r���jsBr�6_�UN't�]�%DV�=��v���Ѓ�[!�������t�/GkMJ�*�&J����5�+¨4H�lT&:��5��<��J�`���À�F��>*+����$��f"�*����劌]� � ����
H�ӏ;�r ^twMQP�����_r�%�f��鬵�˻]7[U�w���ˌф�|�����iڪU�-�}?���K�V�߯v{̙]�価:���Lv��^���c�8h���0]im�ޡL�	����Ѐ��l�|���	�j8\���ĶzM��W���b��G�?G+�(u���{�1��f-��$b@�(n���8 h��S��.��L
K�� ?�9�v�dPɥ>6(޵���K��N}��X P,����?���l ��9Lv����v�ԷhY�^)p��4N0 =*%f)�]����+ioA)���D�_Y��_�	�1���6U�i��'(4d��D��ߚ���D�M*i�e��[�4Q"��c�'Uk�Lz�!��X�Z2���8���O-�K	C�ʳ�/�Q;` � Z��k�B�����&�%��T4����$Ȃ�z�ӛB$냊��:��3���͡�5�\����t����n��D[H�ᏝMX�ɯ�Ɵ)�A%*�Z~�6��O�J+���U�|5)�&��.	�6��M��51i�����9�h׭�ѻ��8�n���q�0f�G����F�@�E���� ߑ�y$���8��96�u��7إxƾm<�H��>�����lo��1tW~ �F�w��Z��6c�]���HA~�F�nDN{������0N�e��>��P���5��ͯ�fh8�bz�x�sI�����%1��Z�`�>r�N�|yV�i��f~����/�c),`����/�1V�yU��O�F��Ct��c�y��7��v�,
�s����P���{��8�q��Er��;ʾ�d
禦��ㆅ�M�fP������z�fw4�1�K�C^)�=
�&];�Ը�k�=�Y=�������&~U	\e�3Љ	�8���	{ѐT6$���wW����|��4aM�.��u�Y���iq�r{�H��;�F(���c�M���;���ެ7hJ�?� ��G"�̌vb�˂0o����6�g�J&]�#&���[�+M21���Y���l�`�_4��:a��>��m���S��x�k��/� �Y���u�����c�H����s��oz��Ku�𨅂����c��X�Y4���j0+O&E��@ʪ�9��
vE��s��q��eb �����FG�����+�>�����_�D���7����v��:.]�F3��Q�:����l֓�Ő��q��мf�*�㌋Z�����	<���!�2�˕�GZ�1Ms�>���Aq�  ���E��e�B��j�}�USJ���0-����0��\�{�*��)ܪ%ٯ�&;�{���՗'o�� #jK��� ,@�b^�+�(�d�4�+��E�C΁*0+]�v/�]ԏ�@p��P�5�ŏ�ƭ��'��b�DY���f޷>b�)�4v户Lz��!��ˎ0��46�����a�V�2\�ݥ��aث�$;�^��>�v`u��O?���m��4��BO�M���1P�qd0�L{�Z��I�vd+2(���j�=�XRSsΫ�R�5��f���6۳�T:*�sB���&^�
E����0����o�f~���lz�2w��gP�������1n'�&Ov�,9�,�B� L�%�KR����M�w����U�T���y\��#6p,��f0̤��d�)#C�����_��d��)��rE�y�ޥ:�R	?�NE��g����) ��>���N��y�����hj٦(}�.��9ֲ���ۈzkL��H����eM\��d߷��D�T��1t-eV ۸9-�>�N��@���߽��Jl�?���L�o����g^�X�A�ܠ�*l�R�U��(v"��E',�cy�F��r����ML�?}V��vrB��Þc���������!J*{�u�/&˨���0�}�x`Ԅ��U��a���� �ҽ���i��D�ZC4���s��>���_�Hh�A��c'�� )?ۨE~s�-W��)G@HLOKf��e|�(O4�� tUC�d7�,}�� ]�m���[[�e�������b"���Fp{���T'�ϲ�2Y������O%��QB1*N�c��~^��[usL�L�2�ɮ^�z�`ǚ$�fpǾ��NiE�,��� T�d�N�}�y �����Ľ�(���'�����KH;����
�;��p�3�:���w&L�s�i'wOZ-b	�-�^��`�]D����<&�L]"�tŝ�*~R>/e?�Iy<��S�33�kO�#_uS�Nj[AS�f���.�T��/GS���D�/Z�M -?��ޫ��N���H̜�\w�'J��	��!�@`���S�(�D��M��V�*LMP�qR����OWNl��ȹ� �1f�REZ��mi���
e�u(��H��~L��.���P�@嶏�9ґ�W���R44S
��o���f�5�����W���~	@љ0��{�;_���j%�d�W'�G5h��2.�\�Wm�#>�|�����dU�m�̟�t�D�l�G�ն�볾�iD�,�_Ȩ�__]��P-���Q���^1���	|�v��.��:�O�5t5�w��$�*�}X��b�8�D�Ⱦ5CW�B��Y�&@A���
է��?L� J�����ή�(6y�K�`�]ߞ�ƔЪnrN�Et��l���[��3�L�#�'�_?�������$�����b���*��yg�Q�$;����o�ݔ)���e��ؒ=�m�y�������]���?�1���2����Eƨ������%���,��Ļn�F!�Orai}���o�!ذ�5�X%��gj$���A�'�WUF�h�s�2L�b7A��.���{���ق<�h������X�8�j\�68'	�u���߫O��*���<g�3Ɇ�#V���S��b�&�,ڕv#�<u֬M�B��Z��'G�m,<�<V�=^hn���ex�F����6���4 �VE�>���aG-V�X���r%��F#wQ���B*�lW��;K��	����Q8��%zQuj1e�6Pg惗--�.�M׏�"9�p猪RNs���^t��b
�xQ�n�6�bF�Þ#����<�0����̰E�V��1��`2��~#�P�i�fط�?I��	�&T���
}�4�\���C������x�i:�
�u��G��)��J�&'�T"�ܲȊ�M�˸�<���[e���ټ�U��a�Fѡ��@�w�Vڂ/����]��^��n�ꆡJb�]�9�`��oW:���Ǚ�B�M�\.΅`$
��<��?u"�2j�5ڔ�D �,^�w�Z��J�IR1wLe������Z��4���Ǚ�J�ΥRв�(=��e�M�V�`"��$l�(Wq`���Q�
��4��(۰�#����;꫞K�A�`�L��Ǭ�mx%�_�otxI
���2�b'ʳ�R���K��M���f�w����hm#�W�����¶P�D�Ϊ�=���`^����_�}�j�=�f�26T;�p�2�-�s.��r�����H��֥�*���K�gw����Nps�Q� ���H��f1��V����ƃ�4<j}���R1���@��\�����+�zJt�'�b���#WeOt[� ׈�$�'�l�Fڦ��*0N����{!�%x������T�aN���"�0�[!D[�Zg��̮��۾�z�N�Nd�*=<��v��5�Z2�k�j@K��x%� +M��)fO��%���Qӥ��K�<F�B��p�ɫ��7f�9�[�O����[�����3\�s���Z3��Bz{�����e-"�݂ۭL��D���_ �f�-���4�һ���R�2��C�]�~�(ip|5��f�t��P�����\�8�!Ƞ��KA�SӐU��F��ޢ��K� jʗy�?�mp'*vnf	�FA�Q���V�uu�~# ��G�^ٖ�=�$����=E_+FJ�]��n�����8�T_`�~	}��(f���������ӕC�q֍����� af�$?�N�e�{���'R�>��:G�>j�t����:�meL!��^��Q�9��'S��.O�dW��Z�����V�n�jl4P^>Ќ��*�g�$JVt�	�L��F�s􅎟]�����VYuR�!�|ĆI�±��P������i
���*�T
+�W�0b�L�;��s<eW-C�(A�2���-i*������T)�np������9ɲ�f&�N[��(B�����\�r��1QŜtܴ�� �@�{NN��l���c/�I��;�?1�h�:�S��n�CpD��*BQ��=bA����g��Z�(��[_~Ih���x��4�{�����
�����0l����L2��WM�M�H��r�����q{9}Pˢ����H'���g�vI8�ȃ�E�O�,����/���ԹW���pk���Zc6���#dF(5�N����6;��J�Ǜ���[��	njL-	[[����Yt���!�6AEA��z��Y�8���F�r�G��@���P��B_OQ�C�|1�L�īw��T�Ц�qiH�t�i��s�]��G�)%� (p���Éɵ��5����lO}�0|��Z����h�h)�	Zx &]?��y��|H,���Q���6q%v{3iq`�������
����9x?�m���wK>�K�T_[��[[������[%���o�'G}vFY��=Tg�q螇�1�]5t��$T��3����#[ɍ����%h�G�=)ΞdN0�5s��ԫ�-�=�gi�v��b�Fuc�n���2��҉[�w��}7Pp�������6���yb�'ƕE�<���Yi��q�o�����Է�4�Us�ƅ�Yt1��|����88�2���>֐gXtz^����5O��;|<���-<E�sM㎫Wg�!(l
���~�] ?l��;r߈��%�2R�x��O���=�P���j��պ�K]G�U���m�fVj���o�r��5�$Mo�bߵ&�Ew���bC�9�4��Y.cbk�~�א�d��,|9^R�k�2�*I�iŹ<z:şYfz��n�Ws�����g`7�T+�?�����T�}��8.�:��H=�4}3��E�g�N-������R�z�~��V>��47`-NP�G�fݨ���!�O �5hR�ܽ��0@~��G�=������|� ��MȼNmB[�!�[�燧��"�\ �9�)���@k�uHq:aC�[V��**�b�zi�+��pm;M�8��H�+�.����>u?�;�u�1�="\��制ɑ�_����9�ЛB5�VG#�k�thZ ��k�bR��,~��3*�~W78���ʲ^����]���L���B�]��Ɓc�� ���]�Uff�ԛF����9}����L��G�[����|a�,���x�'xoIB�q�4f�2��M�k�R�O�M(���z��L�c8��lVR-���1�[�I]o�1��;�w�m����L>3��|�w�R\�j���B)oo�#����8���,�S�oO܃��#{�k�[ŵڝ-t�ʦ�׊�������^�!4�hU�u�H�������U���j�}/��az�|���6�4u���~"�T̼M`�}N?/�穪��Y���w;\��/�Sj�_��ݐ���e)�N;ׁT���� 4 Af�_� ���ud@&�����ƴM䲊Q��d}��n_ʉ�2Ң�r�u}���2��
��!��Q:�9|�	RU[Y���Tb��ߓ����0���v�9t��Orx�a���)f,�m�Q�NndT�'�{M��b�t�׏;�
��[�\�3 /	ma�Sݫ��4�ݟ/���n\�����0��GR���H�rimD} ��<k�I��w%�3�+.�����MH+A@CH�F�S&�%��\�9k���L# x�w;\XTT��b`_!'\|y�B��x�2��pA? ���oR���Y��*�(Ob���"�Rxe/�_x�{|�U��\"80
�����AT��eH4Ӧ�оA��`��G�^xA�ʍ�z�M�rJl�� ����Ur=��D�ꑁH�o�yʾ�e�g}5��W<�Q+�6�O�w[���*�Z��!~��!�u����=Y�z9>�N��z_+G�Pe�ݱVw�4LDȥT]c�J3OvO}|n|]��Cٲ��Sn,�	���P]�XwH�o��,��j.�Db�05���8�r���+3�;��3�˂|�N	��]��ϨV?c�Ο<h��Κ�!�;�E�R#�q��5S����2<�t�N���'�N<���>���y�f��Q7�W��|_�i��B�?�vO���
�y�`l�G
�JK�<��%����	¡4�~�,�c,�d��>��|,�vaEl�|dA(�܋b�!l� /4�̢*ɲ�w߽�����h�&%}��'9�ڎh�q�V�v!=^����ޔ�.S1D���w���VQ$:���
�J�����:�����H�)l��f�?��� �k���ਖ����vTAP�a[m�v��_�ǐ��7���	�7c�9=�录�ȧ�ܕ �b�'X{DV���7~ο�r��ʟߣ�Yؘ��,rf��=�c�\�N�<�#@F����ԟ��)S����%���W���������5������,��(�%(~�����p� 4;]�^aq��Rgq'}	L��v���þ�*���LdAO�c��KE ����J�J���
�O�S:[�����q	��]h-7n�o�1b��?�+]��18'?"c�˞'��p�F_O���!���AȫG�!�����T��`M�
����9�	�6�&[�k���j�F��֙���S �Tj �ʎ��/�p
�R�W�HQ\fp�H��*2�t�Z*�Q�}S�#�M���*�#��f�����q.��5���ΧJ���595$����&Z	�Է�"�5���hͼ��[5��`�^<đ�����3���Y�� 5p��l@�;�44h�IYA�O�� ~�������X�a��@�mx����J84c>̊d���֓'q��"�.�f;�)բ�1n�l6�e� mk�b��?�+������j�dP���bK�ċ�T_P$�i�t%8��Z����ǋU��M��+�̭"E!�x	vĬ!��rШl��^oEp�dx�$��6#�r��I��
f�2�xRYo�鬉�m�v�On�G��׭��Jt(��eF��g�D������n
� |�<���ڃ����M ����۟���mN+
و���N�#��2��I��hu����5:�^���aHYRp�Ȩ;���1-M��c��?&��s�+3�ך;�[������G���:���~x�ɚIr�KNm�K�|�c��FkY�ei�I{B���|�3:@����g���!��'������4|$a|��m/~�BVp�ù]:I����U;�xʹ8��%�L��q�Q�"0���q�Md����=�\���o�T�WC\]os��d���2�W���E�&��ñf�"d�;=��7�K"x�$�x[5G9��'�=u��Ӧ�lꃸ�A��?B�j[2Y7��=]��BQ-�fm'%�zͼk%ivO%����-m.�{��l�1u�1����BU�9$l���*�������ϲ�chc#EE\6U஝��>��|���߮�p3a6�����9�K0�mq���$���"^��<���S?Zo��I�2������	!�e��JNjz7��"_\��qVLbjѢ*&��$Д�m���>�wM��|���v��Kj]M.��T���&��p���h����vZei��@a�d]��H%�[�>�c������!� ��0��dO@��~���g�mu#�9p\v��#p�C��dѦQ	ra KF-/8���ѝ��8�F'��b%B�#��>�ubc�/����Qr���z��t!��3lL/Nq�'v�.�:E���;7�i5�n��Ș>X��Zs��D��vZ�e۹o̊��OqE�s�O�)��9W`�I��ܟ n�'��c�c�b�����Hǈ�z1��J�:n�~��ze�Yލx⇺e���}ظxI��ч����>"��BT�J����(X����H]�|�r1,��k	�^QX)��j_����r���6O����o_�4�}	���`h����\Q������H-�oS/������6c�w:W#��(�FQ�C����!pC,Q�6�j��%�<�'_�����L��C���`c�E\�Վ���T7��Ϯ��
9�E�Е�1v5t����;��.tR�h~Lu,�8&F��#H4ʼ�w�%�7F���]�UTcˡ�{���XJ�� ������n�\n���@�����5FLd��������E0���݌�3��(�J��;1a,��M���}����X���5/�ް�~���z�m�hJO�}�#q��\|���t�y׽~+,��@�&�ɻ"�^ۮ\ !�,plθp�N��K��l�-�Ţf�[�"�M��-��qG}*&az��P�++W�o��U�X�D�H]{h��/�{��O�����X |�"���T���J�4�.���U\7:�d!F�@Rۖ\�-@Q�؛-d�W� �V�{��BDH[�u�������9N`>*YϞ�c���d(�o!�[�K�%6e���g��58�\~ ��m�KL��	Q�!����L�_�*�C+SOk�~���Q[=s�<��p{r�$�d�ţ��unl
kY| B�����u�����I/.�B7�SU��X�a{��v��k���&�Ǆ8�P<|B�\�D�O��]�w��`d�
]��%K��n�m�A�4�2CLd0��kw�M����M��7���>�d�L�A�n�����7�Ά:](���=��{�C��|�܂p�1�!2&U�c��爳�[�����3�_�.P���΄<e�%�D1��v�el֜JZ���n��h���4�8��Ä'�z� T>�bFg�s���[D(vQTj��}�X/��[����<M����9�e�fq@�%���,�~�� viD�72���02����Q��Zh(�YN�=Y�����nm�a@�x�Y1�I�0P�uUY1*4�6�����A�_a��X���P��B��VCOf��k��Mmo����U����%N,�%�����A�#��4|ӯ�|A��M��\� u�����? v��!��a�Y�$Y��VӦ�Iê���˧z�E��]�C �<j�U�/�<vn:�|�㴤/�6k^�o��U������}w޸~�jD1�`q���Y�[�8�u�bmoUC1��+����'���2x\��+V����.U��t�hi̴�%	4�1D{'�vo2	q��4��gxDӖ$�[>J��!T}�qJ7�8�@��Ûű�\{�T�U@HS���7�0~';SLdݯ��k� R{��6��K�IbN8@g,0)6:�td�\S��{�o��IP|Q�4�@���!�F[�cMQb-C	��M5!�<�c`��c��!�8��m�
V�]��n
r�t�[.+��m�����v��=���<�͛�'?�1q�*m�q�	�ZǴ9O���+����#�^eV�j"-'��׺���q���P{��o�b��	ɞzNM� a5 �-��3�e�漋B�Ǆ��^�UMJ?�^��2Rl�q�њ:��;tR£�zoR��<����!��70���Oxre���۰�Ca�L�!:����TZE��N9�zثK� C�~[�A	�v��{"�$<6:�F�>�x[�/ϟ��#81��)`�����pWs��ț3�+�[Gyx���-�Q ���L���)� �{M�5-��
n"�J�4״��&m4[�X�E�lOl������}Z��I��Уq�rD�v��ڋ�#�yRy�<.��0"��ro����A�R�pf믃��x¯��[Y�LW�N�~ETFt>?J��G�	t�*��l�=���[u[�=�[<��0�Fb��[=/y��� ���P]����$�+��:���y㫂�Xc
�)W��	ڇ���d�@~C	hc/��ysAg���Q��b�\�1v-�t��wmK��H^�t_q�@�&����$�P��vq,���_��/���ؓ�u���{��E��Bu~!`^u*�/8�L����܉f��X�<dr���>'�|*�!ְ�S��6)ݰ�4�8�4�����!��^�[Sj0�:h��+%��T�
��[P��� }�����(�>�k���G6ѻg#$�����);D M��%&��>���T�'P�63�~/�*�OSkL<���s�~cp>��\5V*w���̍�+뽏�&q�����l�?�N'	�Ѷ�+`Z�D����>O����9[��� #��j�~��Y���������+ʽ�q�᧱$
�܏�7� �%f�v�!����F�����@a�#]"2Q������s-w:�D�	g=���4�x�#G��\> XU�MI��(��ĩ*Xح���/}>�(��v$Lv4Y�x
n�p��y���L�,��;�3|P�־����z�x8��_��8��!n�B1;��2���`Ѓ�%�����A*)y���'A�%�~�^��j7d��^G@h���H_�2��0ܹ���j�8�"�b���a�8(�R�;΢��iQ�<��z�b̯c7���]c ʤ���9 ��� ���}�p�2�1H
�.������D�W|w�+Q�Hqp��͜^�)��`�${�'��p��7ef�U<0�5ror-?+���cu�1�Lni��(1�d���a�x$|gP���|�ku����~�!X�J��~*��gcF`us���l���;,��-�Û���iLoq��3
iT��B�F}04'c��:�l�E���nкLI�:p4�6: ��xbf��@F�θ��;OMF�Q8��.����*�0�8l0�Ɋ�����D�=�3������^�R�aGb�X>����ڐo�@丐<�y	���T���Xx?�T{"��=��b�>$֜e��"���x׎g�l�A^��jZ�*�Q&��	:�|���T���-"h�]y��;��sS���a�y^�!�-!k��ꩈe�=��\e��d��dV�~y�zR�H��D
!!��J>�|��aȇ!�*!����x�]�������"L>�	���� �o��Sf�Ni����V.�hu�������J�+ �Y�+8�{��-�a�DNK���&a�gcL�~ٿ�̄�q���{��"D���kD���X�����>�!~.�M���'w����\^}b2m�l�bX^w��OG0=���U��1C"5=j�!�;�U�p�b,>��1���[a[���b��T�Z�tk��P�Y&�ط@cf��`Cʞ��sأ!_�:fA��65~9�k�U���|��܀�*܌�͔L���5���Pg��y����j�_�����]x_��~ß�2w������0���b���&\�F��:���5r�c,GMM��Ƌ�
뺐3�e��5�G��c�r��Xi����i��
^���bb�G�R	 э��,���}S��ÀكO��~�Wi[��v���b��eJu��A�m
��3=iS�5~��ߕҋ�S�q�.�Rj�g	��j;Q�k�!;�[^/.�w�hnpͲ��[K��'�o�
�dQ�l}���~2�5(�h�2W�ث�˦4.�������=?��z��~}�;aL��D��h�0@��У�v͢I���7��Hu��j�?�A�_��T�����.�#�]�V�@�I�*�F�^���nd3�{Z�Z<^P����H���חV%}I�˖X6<t=����vׂ�C��N
V�jUư�?P1FY����%]Vtפ�=���<3���9A}n���ڬ��i���6��A����e@��ڎ�B�'ԛ�4/MlA�g}bݜar
���>#YJc��N�ƪ�||�	�FH`����
�eF���I߷�6�o�L2��M�p=��MS�ڌ�=�sH,��Y��{����;�9���P�9��g��@�A��0�¨r{%w	.Y>l�/�z�U��{3C��T��U�Gh8vl��nz�-�����!T��w5�6I��Wڦ�ƞ��z6�Cݿ��%xS>���sM^ڣ�;E� O+�z9�KW����M8�h�@,pV��W 4:���-��O-㢟�u9�.2������V����H�>����}� �Y&�+�m�C�^/Ի�hZ�鏡���:�mC���|.�#��zΙΤ�j�K��gN��p]/IqfAX�W4�����?�ׁ����Cǻ(�޷�J���M�'��T���"Ǣ���DOي-�]�Y-QQև0"'�47��p�hʬ��AƯ¿/�������2�zx������������U�T�.$�6˶��S*ۿ�6D����y���3.#�;cf� �Aʋ}����W���JP.8˓.���V�(�E?ng��-��+��G�;�j�J��RWe���
N;pP5�.������!e�C���3�7g��gg�m�O�6����SP�6��0�={`��1CI5�����ǣ�a6_��q�/��;saC�2��qܣ�,&���(��F6��gH3����:}u�б�Pb*Y�"�be��=�����}��X�S~].S��,K`�bd����П�"��Ag4Y���50D�[l������;����{�ӐD�(=����j��df`��-��lQ�Ԭ�<g�9ҢU����{��?Ot��m&������;2.%y�퓔Ǩb�W�r���*0U:���߇�dQ��B�r}��Lm?e���Eɏ�#%�^��!����H�},���6ȰXh7��������e�_98~}VO���W	��o7B�O�(�W�s�F���1`�``�P���bb^�X��1��D�����p̽+&��LbK��&�B>��=�RK���$�:��q�4vI�E�@��^ aY�%��n�n˝�Hڏ㮻�)rW#n���9�U�{�d�踕�,VZ���d�Χ��U�l}|B��/��:�	�e�S�H���Q�*�+��߀82x�(Ыe.Z��W��&7l}������IG��,6��(�.1i@�06��	n1�O`��ϒor��J~��p&݌'���~:�����7(�(Rb#����7��R��!D�~jS�=b�
��u�H���O'�z4JP�p�]�T�!����7�tmJ)����BXZJ�ъHH{�Ɍ@3ܾ�빞�� &�ѽ�A�3�aK�?�)�_lZ���E���l�$�p���	�n��>���% �^M�Nx�'�c&A.�=X�7 V�a2)Ņ���٬4tr�-.�De?6M��1U^_n��  ����'dK�����Wd�8����%�"r�z���`z7N���[��V6O#N���X /�T���-�ez^M���Q��������Qz�':�*�e���Ja�����Y��猬;�X��#�DL�G�4P��.#�_�7ojj�&_�M�N���v����uv�g����>L���D:+e�:H��F�ՙgY�,�L,2i�Q�d���=-*O����N++1��@ �~��DaGA(��2AP(HW[� Z��f{�<�������(
��-��O��#8���Cy�TJ�wp�3���\�{(���M�Sl �`�O����VUư��aS9�y��.�:�PRʪ��e_Z����wE�������#�����^?����/:�������,L{]����d���"�h�?z�E����%ߕ�dD�W�~)�9��c������%��*��!V��g#7+4I�����~�+�3i��p>���#�F��.������>y�aq�����MG~cR[�&ju��o9�s��-!��F(�}}Ϯ�y_nb�|=�8ߍX9|+^�ӥ�=���~�݋Phʜ��A@H��Ov^|���=J��i�^�s�$s��z�i��h�]þh���n��f�İ|�R$�(<% ��#I��_j��y�,՟!����8[WYK��x����*a�� �0�ٹ9�p��H�x?C$E����Q�"k/��K��z����;�e OViF�~���K�0�r�<{[I�]e�`��s.��ى|\�r���5�����&��K����,"����צmQ����Iχ��A��L��lA��Y9!��w�h���냵�.t�n���6]	�q�ΐ;���pZ֊�)Q���ԍ�m�T�>6��+�U�w�Yv�A�o�5�}+���ј�7�����P�M|M���ty�Uq$��!ۣ^2&�R��>Q������M�Z�'�D��'ZH ?٘]�6�����R D>�"����e�#C
�H��}����*��Ú��5�\@�"�5�m3��'M�*�OI$e()J�)����)�l��A��Pw���m������C�Zn����a�+��J���a����p�����M�B����Ά`�X��ҟ$�<�d�_a��ui⠚���d������#<�J�4���I�>^����) Ζ5 �����V����#�;+���8�>/u�/8�F�x���B�C7�q��n�bt8�GSRT���폷�u�h�Te�z��S1�i {�T	2�2�|Љ�N�5�8Vy�ލjT�|�����FV֦���@,��B)�]l�s4�3�fR�="�&�������H��E���{\�qN��ަ)u�3����7�.��<��r俯E`^)^���R���?�1���R��r���	r41��rz��D$���0z�	r��ߨ����:�3�0��T���;�=�3vq�4?o+�0�.+ �yƇ����@ߥ�3:|@�Y��μCt��ܤ̋
��ט=f�8��E���m~`�m����+��a���zW@o�D�b�_��h/k @�<9-��rT���W��;$l>Iѭc�uJ���t5�?.㟝�9���t[6������x�O >͈~[W��`a���"3E+�T~�?�4U��c�� V��ZU�s"�~���?��9�O�9��mC�7�JI�ʰ�U���xV�f�d�H�q�l5̴�qR�X�0 �����i,�0�Z�,I�b�<�T��r�A��ď������f" �}��5�+����^L��~�����n#2�|p/�l�q��+6%��#�{X�gn�H�9���\&ݠ��H�w������y�=�G����l3�SU��Oc��)P�PL:��pw��A�(�h�����g�i�f�`Q���b���
�U��#+b �bm�� ��|�� Q���R�&��
qE�̾}�����Γ>{�A�'zbB�:Fb�Nj��N�����j�����������1���	c;��$I�K>��x��z.2|Ċ��ґ:߂���qA� A�4P���9�ok���z���x�I�w������	�8��x@���W/�я�I�;Q���p�f�H�X5�Lℇ��R�����}Id�pA/jqci�|*t�00{�l�ӂM$�̴���x�97�4g����[k�t���i�<�!�����	%['����f�Y�S:�q�xd��a�����H�F�Y�'�x�-�b1��m��l�@�~���D6SbD�&7����H�Q��i@;�D�P�8��7���ژ$j՟��[?Sg<N}&敩Yz�X���G��e9�-���-�_m]�F��$�Ӎ��:\����{��ij��U:�?
6�\��S�.d�?[�����n�t�j|�t��ؠ��������*�#z����0��t�{��=g��lr��Q��I�H]�*�S��h}\7&_�],	ү鈺��e��]�,�@�9��4�m7D��;��J����m�o\�ڒPtdv����T8%t��ܙA9/A���S?9�XoH.c��Jq2��v�̕?���gΖ�'�(�=�1�&����E���|2L�C����^���(�_��u��e����%�#Z�7�C~�g�~&�B�Z��5%�C�`o���m��	���.$�):~�}��SM����2,��ڿY�ꋭg�P;n�� �)�E� G�&XE�~\��}�$3���R�<}�����f�F��<>��n�~�ι`2�S���pn(��*�O����T���f�G��+1�*B�:�a�!�/����RI�YM��Dq���6u�gxo����]��1U���>�q���/�����]�p�?5>�I?9P dx��'�{q�̈́�w�A���pg�-9���/�Q���Cp�g�^�1$�#��q"�`;Mk%b���M�w�⇘�������W �����ޜ�&�~ʏ\Tsp�e�4d'�տ������ʡ]Z޴���ֈ����FQ}����@K��Z<��F�E�G$X�1���N��D�W4���x�ϲ;�/Y8�̾�&A�ƫ��lvo�TA�]�Ӎ���ӳ��9y�b����M��ʅ�����ݥ}N���d+�&�qw͝MXl��ё7���FI���d�0�"�d��
����K�M��p�&�N�S���b�H���œ2ΕQ>[�O����ũVwp4��UוTߩ&!���+݉L��r���;�'�I�S��e�㢾)@�B[ ��ݾ�[���� Y���u�����x��p(� �q���&�,Cz�f�-0>���Ip�&�V~�+�B�fP���fC/7<o��HO�t����v"�GpR�y������x;�����q8Ǉ�i�E��������Ʈ����<
 �PP��	.�G��֨��.X
7N�vݳ#/ֳ��H�%HÞ�8'�����|G	%\S��\�"��W���,yx�:���� ��Kֿ��%<)�X��y+�EpFu��]�C��&g	�8�m��(��2>���X�h��k����b��q�F�j�����`��œ�������z�v$�P��7��.���F��F}ؑR7\�\7�lm�<V�+6�|������!���\�~DU�$xyo�?ZuF�_L]wR����RY�E)�3NC��QC�Aq
�û�9S�J6���k�A]މ��uo�P�]�a&.r^��Fr��P��d���j��Cs�C~Ы��r<3�nè�I��hv�7�Jfb1���Ď/������E@y�z�_2W�d
\��T�P�q�獺��o;�;!�ȕ���Y�}���qL �PX~��G��wPǵL��!��ڞ�����S��"I����'>�ol\jѠ�(٘t�x���j�ϯⴝ���� !K�4��l$_����%ɨ�K���tG�'�� ��*�׶�iv��W�����=����A>�*Pe�/2u����Q�I�S��<�P���}��K^:�o�\ma������.�z��@iI_��������ׂ�<�gw�wތ��\%��G��]5�۹�t���
�Ҁ{��8�J�����N��8/� iI�v���"�,�m/c��3�+9˗�$3�0u|wA�A�}󽞑O�
Hm#7gW��j 6g`a)�Z=��-��gUA�򁎦���~�[�P�/y� [�T|` n`x���1J�[|p඙x6�P*z�쑒i��[��S�G�mk���C��j�!�0j�"my�Q�R孏���j;`Ƭ�2��ĉ�!�S����7�-Q�,z���@�I6�{ o�>�wP�K6̸�͘8�W�_-\9����u�^D�����ח�ޞ�Sdђ�{����<���L3!��� � ��Jhg�xt_3ɛ��Bb�(I��?0�>o
�55�4prČ?F�WA@e�D���4�Z�´��>Ռ�x�#�4?�<V.���������h�qr.�P����u�� �\��xb��ڲ� �("��Dc=��Xz'�ֈX�{W��տ�O��i3��4�aI���y,��/�´�4��@4T�9��X�Jz���P�����%h�)ͨO�D����O�r]�^B���ä�K�|�%6l�EX�r�Y+VTy�f:@o��Z��x:��
�,1-���������]-���1�&D5�@-#��GΪ�>��*;��R��y�L���8����/0����b��N�^y�=�,���Lx��l��J}��+�	�C]m���Oc�8x����/�_��p��J������}F��;0T�a�ӫ"�6?nn���h�R�[ɫ����ӛ���
�u�)ї�8�U�;KzT�Ac�[��|y ��5��a`fIRn�M^�*����#o��s�?���]���)�v��w�G&k������R���i�6��R�#:�@�e��3(�vW��)���GV�t%���i��:�~>�D�t����$��)�FC���Հ���gD&@S�Ac�%��'��=E��K�!��)�3#|xk�����<}@�]��gc~�Z�IiB�w�)��;����qr�����}	>��� \M5n��/t� �I�)>��e��bB��Y��Ձ<�f[qN-���Z4��Wz)Y :5B'�߆=7�>o^��.$$)]��`9P��aj�@���Q�F��j��tgդ4�\z��G���<�6�,�'�%]s�1*]�N����H����>�gh��c��9�[�?�ɳ�s�|QZ�L&�q���em�P���r2�hZ5�+2��U���s����Ј	I���p�[�%'z�eG����u�S[��fg%~x �
xg��g�������s/x��h�v���&ݤ_�����$�<��{ f5��p���-g����!n��Dc���b�G��Fp��c��{�Y��J�C�)� �0�[�e��3W�Q��(r�*��{���5��7��n��z�MY���b6��YZ�|�w�m)?�NU�����(xq6�+�׋W~�m\�1��+g�'ؚE�f�T[kD0�V���&d0�r�+ڤ�=�Ex��g	�R�%�2B�y�W����l-�\��aT5�0&�eHb\��s��e��9;���ӌ����ږMn���P�nU!�o����]2k�r�.�i�����[u/%�p��x�O�U��e�.��>��C��F6��^ �9 �����TDJtV�O���:E�(�9Q�2��o��-�Pwd��S�XU9�Sw:-���I^��φٷCŋ A^�!�p���j[��&
���8_����5�IP\���% Y�k�<������n�r��e��v�}=���y��_RoN��>G��? A/�v�
����X߳�b�:<	E�I��mz}�wM�u��B:��it� k�*�q�)xlh�b���yi���y������%�ϣK&�!Y@��o���0\ρ���˅�ސ���k���r]�(l�{�\)
A���g(c1���T�R���lr��|��!|�_��"�v��)���K�,4��	���Z�:�ӽX�LF������Y�LR�����igt�F��&��j,%k���2�����)��ۃ'��K�L�����E�Lh�&��w�'��#�NQߴ��41+J�&A��rȃ�`� �	QU�kJ��0R�x�U�%�;�hdE"���ޖu�1�����a`l;�m|fr	_.cW4�Ñ�0���A@�a����&���¸�,c*�D{۹i��D±�<�ނ�\X#���:ZE��C�X�l�1�x��w~�>_�
m1w1T��)���̫�x�5r���k�<"R����G%@��Пߠ*9ᒁ5V��aX˜�qܜ8���~^J`z�(��YA ��U�ke��w]��2��	REG��,'MCw,^�G���q�bt�}�&������(%5��qk�6"��7�В����#��
E�\�9�i�.�0fI
o(�u/��w���M�Vkx3�^��	K��#��*���X͔I����n�g�BU��0�kp��C~�
�P� $�#Ū�u�����^���O1�3�g�?*���)�Ӫ�]D�w^6�^^96.�$�����k�=>��㡼�\�Y��{}��b�]ij'M���f9i�����6$�o%�s­B�m|}�i��-��j��df{��dhEkiHA��#�cw1��5�_��o\KNr���d�˃%�ߛ;ۨ'��p�-`�(i)D�m��Ym�y$>P��� ���VW;	w5tVӇA���,'�4J�=�3�7�Y+�Y�x��ȅ�ԟ9��rv���Bu�ܘ�.��@%��Y>�Q������fԗ�>������	'z�S�^�zך�C^ت��a��待_�g��ě��Rj{�������F8σ�nm^,��`�����uYɓ�V�	�ccN�V9��p��Y��=�p��.�7UCdø�6�PFtدWl�zN�ƒߏ����R�� �qP)5Yv\u�7Г#���,�,�7~�IN`F���5,�z�R�"��9��@��s���<��\f�Y�1m�9g�FT/����6�ER� J�p�<J�u�jk�a�CK	Uh6��'n���A���7qa@r�
"��4SQY K?�/��;h���Ԙ|��1������<�*v�#Da���01A��3�̞���Hp�<��\��h��Y!ۋ��@=XG�P�MĴ��P�a�lM�E�]�%���_p�z��d�
�c���L���E�o�Us������le���ؘY����!�;�,}�D�����||������
�|,6q�r�:�s���	Q��^�ɺ����Sp���w����`}����.4qZ���aS�18�/t &V �����}dǰ-��|^_��,W˝TL��8MB.3�:�(
�K2�3���E��8X���(�u�%b��1W�2��3%�;5{}��z���1/����*-��G��b�v�/Hݧ��6��3�u��Q˳4��9 �g��Ưꖝ���X���A�K.X��I��a&�?��_89n��|Ɂ(x9�RJ��\���#�<F�	G�;]de���_E|t7z��i�֊k��`��t�q���OG�E,�>�)�.�|*a7`���g_J&�I�{��3?�KΑ��� ,���_qv��ې/
�����ӭ�M�����w��Fq�k�:����v豫�^N��NPz�����,B"В�}>�U:��g����و�j1��\���u̒�g5��-��|��J�V�_�#�)��g��6)[�6�ja6�q��dRg[1� ��������2��Ez�8:�H%q��%Z4�3�H߃ �"�J���9��B��ޢ�*���#q3㣛m�����2GD�� {��Ƅ�U	�,��I�H�p�G�u�����#�%Uj���1p�j�]�9�ũW6���_�����G�٩�A��Y����%:c��pb���9����1�4�/J�f�*&c- y4n'���}W�����SV�Z95��(�Mdoa��l3o9��4UU܅m��md���5U��eP��x|2�i��b��R��K�L&�g���P(�4%νL�@S�Z>��[�7��:�'0`��'�r�Pn�톗:�74o����E���&�W-�����5w(���`5��&�O9��" ��CU�  ��BrS���p՝�^#]�vjy����k�����GZ�l���e<��[4q��0{��5�'�^ʢ�m�.�gX�%��䙄�|#���E��ivT�$:;��a���7	Y��2�����,|�Es�n�O)��H�O����L+���;��+yQ��h����u:�p�҈��$��H��[r4џ�	�v�~��H�U0��"�e�7��K�,��8,�Df�(�!�]���C���q���B���+▢�T(k���K�hڕg��{V=jKB}%2���'�N�.����Z�Ţ����s��X,�BS�	��f��:.�i��V�8L�M�2;��<��hYN��Oq[6�7f+�^�̘Q�8�v��Z}���VH
V��`Ŗ8L���"�D�}L����b�k��P5���T�\�AWZ���q�瞧e�;�w��Y�CI�B�Dsd얚?��Iˉ��y���6g�I(��#�ڿ�����	N'���C�%���a12_@�m�!{�`�4 JS��!�0kx���m����x�?]`J֬�0
�6�e�4^Q�D9W=�����>W	�q3	6f�
�$N��􄘇E,m�P��D�n��jɦWPw�s��±���U>՝���k��젞⿑G��,���&��A�.h֙�A9I�w�R�SL�" %�M9M�L5�C�E���t���r%KNf�h���j[u��E� �5�`���k��︋��l�3��VF~ܨ°�=:q*)ã��${��Ia=�A*J����\X��S�#4����_�^�t��b�>��d���ulhs�C�t�?�Mp��k��ܣR<g����I�	�iQ�E�\�g��0��0�qw@�-�3�֮3l���K$U��/vG$��փ��O�=�f��\PEUHñB�G�c�&?\�D��3��81(��L�a�Z�Z��Zj_wᡶQ�pi2[�cz�_d#�"R���C{��$>��#w�� ��3��L�V�=����RF3ZX�ʩ��j���0C����>b��5��xe�Se p�b���2U}���!��0�b��@ȸ�֢�*Fa��*�#�����AI֟���<� 0D�@;VR��éh=�z�4��n"�d�>|�X*~�����56�9*���)�G<�R��\���dۅ�y|��'�m:+�g`E��Xn/./�,_��h&����~Zߡ����}@Q��M0W��������?�c&��W0RB�=��^����Lg5P����O}-���;��#��4]9t�H,�ԗ��)�k&�����7�)+2�a����$?���\�b ���Oh�x"H�E��K���$v���`)Cm�3mW~, �FT��-U�3���h��K�`gR;�n�p�:�4!��o�T��v}FQSu���a������C�� n-0Ħ�3)L�5���1�����W%�+�/>"I=��eBԼ�k|��T���L]�^Ko/O)#4cv_�?��~�\�k#��IT�*k��s�_������bq�l�LZ�d~q;�S����<g?�Wy:��A�U��a<�԰�/�
ȝ��0v�:�Ze������:�4i�2D�4+B�'�?����v?2���:�Q⢇��)5� ��u� Z.6}q�l\��t��5#ϩh6���C�u*�uE{e��OL3$�]�vAp_h������3q��l��;��<ŤG�o;�������?��
��u�_�%_����Z�.�,�L��gܞ&|�t�;��Y����s�ܰBA��?S��[Ǐ���4�6�bSH֮��bd5}�!J�������")��i�20+m"}��X#��X���5�Q*�!�JD�k��������¿nӹ:B��|�BaU�7�Mj��kt3g;�܍�����nB����0&mpI;��[����h�@��d��!u�����m��I��+��b�����gM��Dj�p+���t�Eǯ���n��N���,�A�kW����ޛ��p	�|qh+�>�E�w�F'�9�Q�r�&�Z���i�@����s:!�ʍ�_c����.Ի�t��&du �Fm��$?6��0(y���%��r�]���W1By�����S�������y�h�t>�����+"�	d�B"\;���q��T)�.T��23O'E?��d�gɦ�t�J+��'v����j���:�5��_�:��n-T���%���6gTJ����'�t�0q��1n��R/������h�@oc�����~xvb����}�!��dl�E�>��*�s�8x�������e-�	U�}��Z��!p��� xQW(��4�L��]$����K�?���atn�ʥܤ���\R��D�σ�J��ZQd�T���;���_���yx����蓦s�siq6,�!8E/5_d5D�#�ŰDY���BlobюʜxZҸ�w��^�@�A5z(>���kz�4H��C�Ps��3�O?�	�~��{-���<��a�#&���ۯ���D�HL� xu%���	� (�(n��wCC�"�2� ��(���F/��e�F���&�ˇ�Z��(
����A1Q���򛏈�n+*��A��hق듆h�^.E%H�
�9�"%#]�_H�<-%H"	u%m)�7o�#�!�������9��+�� ��G�,)0r�M�m$O6� K�'Q���w�_�tm�B���qơ�޹�n
"l�֑S�� I�'��ts��}ƚ�1Vk0"�%l����|�&QZy�����;��}�Hː���|}1��m�d勮����^�_���~
�u�S��$��{؛;��t���LyA^YZ��jS�_f��0Y��+T"�FJKa�-��m��n���&F��*�a>]{y��!�,���$���W��	��[,"���H�0�� ���i�,)؂[�$N��)}�<$������`�����16�a���%�N7x���=/��͕R�=י�
'�z�Ozi���^�FA	!������!(>���"� R�,�R��;z`�����^�n;zK~�s�z��V��aDm�1gk��	����Xהm��mt����Er�dy�4�.7$IjȞ���,J��r��Y�G\�̿x�Z'm����P�ۏ�BY�M@�=Z�^%�8�I�:�.�V#���,,�mO��;g��M��������W��!ޱP���dB��M�����z�)^A/���=�5�Z��
6���~)U��Hh����#��`����@XO@�}�U�W���/Į�����wg�*g(-'\�+����2-B1�`.P\�.�� ��U;��r��t�g��ou����`rODn�䆂�z+���QP���̍�z^��|���Yp�O�>�K��T�&��'�'x�T�]EKz��Δ��N/@�O�wt=����"�qdzj��D���vl21L�'G��[����{(��N@3��y�O��γ�T
�e������Ņ�L��sj D(:��5B�w0X��fi��)ņX3�����kX�Xmɒ�d���uQ����^���ڹ�]�T�ԁC��I�A�l� rX%�%� �siqnv㛪�}�Ӡcǘ�1)X_�r]�wT{�0�&<�+��%�3�!����*���c%8���-�LB2�6��J�HJ?OB�:��h�Ġ6<lw-�ԧ��#e���s��	,:W4�0�b����:�t������LT���AC>�g�l��r&�,�v b/��E�?��'�i-�bA{x�#?�i�$ħ�/��4Y��i�:�SN���(N	���P>j)�����/���Cc��@�O�����$�CX+�*|��j�[���?Vm֦��Z~�K)�/��)u�>�W�a�l"�)��ѡKg�J�yV����pt�հ�J(�-t��R�
�bIh�L]�p�z�>�X�����:,����(���<�0����i����|�GD���(��%���ӌ�����w��r�ܓ��.T"GƟ�B�D�Z�э�)Z�.�?�킶��g��ӺnquC��:0�b��cd	�a��%"�L;H�M��5 uf��ٮ���LrȇsX⑛lk*��!��h�2��éY�?�V�Ҁ�Z��u���&�����mʤ8��
ig�"�r/��R"ñ5�>i(�H���:�ﰓ!�0���V�,��Q�AU��pF��k�5-j�gmݱ���H~���_0���9��O��G�/�l"%-�t+�ƚ��"�qPu%*��'�b����jKz�@��#B�7$�����U$[Y�7)O=�,�J���%�܋"�q�x��S���c���KV5��P/u�c�q�[� �.!z?!��T�k[R�$��p� *�-���������Ezs�i�$57F!&�oxH�d�*RVu4��M8��D:�č��eJ�ڂ$>�
R�񊳸��PDK����Q�vt3�%LK� �S�Vɣ�&��[e�W�u}�����	5K��H����(?;9�HA����>���Hy��I|e�;�.Y����jgm��C,)^��1��uwE��e�1����ɎMH�ԣ��і�1��R����aLN��S� '��T��C*���̒0Z=!�P��?��9���M����0g���̑cկ�YD�Py�sՕ�纠�`Y5؋;�뽕>}�pǲ���dJ#�~1�a�,xKs~�BI�wV�0�%[VT�`k����L�J,�O4I��������U�ё����W@aW����T t���JN�Ĵ!SJ���e"$S��&���+p3+<?�J� ��=�h&����F
�m��Ծ�A�Z�,
^j�5"��כJҷÌ,�:"����Pf��
����j2V��Ll,tK/����N��7����}��#���`��:/��*(9��D6�%F���6?V�e��â�\�]���{�WA�����m{��#�l[�Q����}+ƾTQ�HvMJ>Tef~��	�ޑ��D����0
��Yb�rB��W���TՋ�I�"Yۀ4o�|����iQ8�=��K�{Ɉ�Wќ��(a�W�?���0NHb�*��0�&__w���=�E��� 3�����eؓV���"vk�U9���H`�0:��f1G�nZ�Q��C
Ve��8#���ρV��Ҿc�U<x���&�/n�������}0f��}�D��=� �. �h��͔�u��h�ӫ^�z&���t���N����6��d=�]�0����=>��i�e�׶1袧\��"��F���8|��34��?AA��=$91��>L�`E�h��$ ��$15EX�W�gŞܧW�������S�"3��=�Ņ�GRh	������d������fjV��+����d���[w��h&�-.;d�S4S��Ԋ�$U'Cyh*�D�(PiN�GQ�����$n�ʞ����8�L������'�U-{�2"Ø}}Ӌ��橧E�ER��f�Z���Ȳ O8d;�C�\@:�hі�/���S7}���Pk
��O6S����N~a���%�p���P.c��_hI/�w���ˎ�r���}���-z-W��1�L��qJ��L�����x���tu[N��U&� �zR$&��n_������#������O�m�Ӌ����[%Q�I�F�o[�B�9�3�Ǹ*O#\]E�HJp�(yў-�'<�<���#
�����W�vL�ͩ/ ���YY�;���C>;��������-\��:r1z����Z:|��c=,��F�y��tR���6����*A>Y�AE롯6GE�/i��f-������JZ���!����Z0�)o�z�2UG��_zN@� �-/N�p<x�8��j�Bhy��?�3w�y�XX''��9_� �$P|y��/Y����{N���A�mK���B�RGmʕ=�����x�d�q ���� ��wY6Qܪߧ1�-���)��[ ��/?�;&9��Sb����*B���
��U�X���q�Ly�����{7kМ�%L#��ӺxR�~�N�%�J(�	��������i��f{�K�Xu
�\�)l��%j�������p4����`�-�<��>�19����#���_	l���&L��k����f'!�$JK�|�v8�E�U#�s��OR3��}$g��  �6d�v�I�߇��\��ه`�n^��O�1�`��<+$8[I�bt1U:��$��#��;���LS��;�q�i�(|.� fry��m��wn$�ev/�(P�Fh�Sc$�qFo�-t��F�ߜ'�����d��
2>�TQ��s �SXy
�m���f���)V�n�E7�p��6���5oCz4[��]��0��n=m�]�M3z&�������i����t*�m`�,���B,�5�%���r��GN��%,xS�Kį�6�>�z;TLǂc{� ��ܔC�:\��X��jK�?��v�IE%�d�j�A�lSC��`-����E�m
�Go�N-]�����뒁W!�+�}�ũ9��0�R�B����>ɠ޼��\���{˹5��1�\�×��D���R��o����R:f�	�i���_���	�SE���(�:^���v�ȩAH��>I�o�N�SX,�m9���+�/�0O&���A��6�U75��)%������`�k;����a� �H4$&�$'9A��{�$3���*���Y�H�I�	�U�V�i5 Cm%�UtM����`�9fTV����u�CvB�VI�����S�"�iЉF������K/��ݪ��G��:�HyK�n�a�p���q�S�x�<C��ͯc�Sl̗��h�5�?u�ڨ��e/�+F�H5���R3e)m 5ON��HT��(�8��$9	Dg�����W��
�9��կ�j/W����V������9�l��5�[ǫ`{GpTϽ�dP��A�uo^i��y��?���X#�)�_L�nf�s�x(ck�	��괩9�!�W}�~�JY�
А�)�P��
��=N ���o�����OP�>��X�y��V͝�rc
�B㛹!�5!�A��f� ��?�H��H�\�R*����-������pZg��m�U���b���N��ƣ�Ph�RC1S��^	�y2H��7�tJ��5��4�.�S�ڇw�x�.��9��H$��Y�DⷺH��Np �m9j6B���)�wm�9t�|�b��R�amy�t��&����y���3:n֦D��n���8�J}3��u2���Z��;����f �1�+���]�����낛��#�I�T��3yŐQ9vAN���'��q]I�1�w�)����- /Y8��AJ�esa:^���3$��i�e�����I�9�
����1�����${&b�t�Q���z�֫��%B�G�ǅ0$��8�F���{z
v>�3�Ps ��tR����|`)�!����J�����<þ~��7���ź���
��/�?/��4+�=<�8f�B}����Ch�@P�0��p�{��{�c57W��ŵ�R �P)��A'��!�V�i#�r����/9��C��&y�g�d4R�z}���Y��"�S�yG:)��nq/�n]�$5�b&��x;�a�|��������/嚧���]h�%��Iv�hu��D�"kG����|.���*G�>�UYFX�U�F(��4+qz���;�w�p���];(�VL,~t~�͋T�t��"h+Yl̹0@��YI�q�,�ϣ���׸o���8q�ѵ&$R;�z�=utJ]%;�&/��Y-��l�A�Jm�VZ6�y���N���7�C�ʒ'�N
Yg
�%XXF0��V�#����x)$6����R^�5鵭�ٓn�fnξ��)�0t�E����,���������x��:�ү��(G���(K���7��5Ɍoػ	P�z�Ii�Oe��q;n��+1��Z�K5U�Lr�w�WƩ�"r����a���d����)�"�u�`�:����`��A'�G�\�J�-��g��Hb��D�t #j���7�i���Ñ|<#-I�����q�S�<�?�9��Ԇ$3�G�6��b��Q~�N�� ���;q���^;������L8P�������F��F���҂�&) ��M��|����ѥ"]����_�8Fa��?@ҡ������Ň2�	N��   ;o���t�4��C.R�㋊�M�R�%�%�dT�W�>"~$�B<��9G&Ni�Ն�2�KoX�TH>\)�4ߎ�����ރ.f���y�A�N�N����J�}�G~	�=�"'��ܒd`O�Ͼdn9����-�w��n�ddw��ηo�2���0e����7>���������T��4�O?$� ����&#,*V(B48x�_K��nk�"0➲����Pg��P�����U���-�pJ
�v\ň/Ha�R�s'\��J|C��/������[+��Y4��W�X�Γ�e�_g�0�~ۉ��� �ͧ�I��V�sP�0�#3J���|��숔i���c`�W#���z�;`��m.kI:���{�ln�.)��k�����)5�3B��_�0Mm1�u2�%@��{0�o*���W�ۂ(.�1�܆�9M?	������I(��~��3"�zP�,��
a���U��� {��J���:	C0rn� "�u��Uws����! I��æ��sIF������� ����
���^��t]t�7�(�`��z)C��J\`����Z?�z�F ��I?)�?o��,/�b�p� r�ex1.�^E�t!O�>�Pfº���	GB�-f�UAwg\F�V�ca튷��z>����graH�{��¾��^���ݤ�!"łd��m^YZL����~��k�v�D���&l^Kۺ���R��.6�U�b��`q�7��E��'*�s�Ѡi]%K���}jUtfqR$���S��#����'� %@���D&�,���ð_=����YP��X�^�|#%I�Y�M���Ƞ=pfpfD �R�|�����N���bm����;G�_خ
<�%��=���P�����1I�R^��Rq��I8����ߊ[]�n/dw�����,i��w�4	��J#[�"�:��\_=�ń�?�V3��g��M�R����"�,f��kaCm��Mh�f'�O�7}�_,Zj�)F��P�`�F�w.V�ٚ��ĕq��a����W�3�>��PD;(չ%���Z�g8N��������%@V�Q�9�&�������-���YK�pE��~=z�W�r�%L������t�Cy?�<�+�g/F��[W�O6ݛ��4>���b�h3v�X�&LG�xd�.+l���`�v$�b2�%ݺ;��HU��J��=�x�t�)�"�&gԢ�O*Շ��y
U`�y�Ǆ����W]3��Y��dy��X���B��ݎ<Niy̗cZ���QS�u�f(��Q�����;����&^B���,_�`3ÚXǖ�Tp8tW�Ah�F����&��?!$�,G�D�Ptz���2���E���%�~s7�I�Z;)���vM"��<q�c{?�����T���R��8��yĘ��2$��4�&"�D,v��ͯ[�]����UPqC�i�uȸ�Ɔ<���
�r��.�]ZZ�@U�� |��$O^~
���������x�c��e˚Z}��%�	I~Qچ.��%�y8l�� �x����sa��ϓ���s��n�KK�쇌��R'��3����٢=�	����.�@��"7r�U�x�5��7?edϢ2Q���tǚ4�N��:�2���Z��;����LE�����BUvF\,4 ��$I�[D�����LQ�DNp��{�֙j��YkN*�bA�ݫ��<îw4|�}a��'Q�����X�taR���V�����v�	q�y8Zs��y�"��-�ݓWP
s
���vxrB3X�=�aЄDY�aC�	�#�ЎX����P��F>�b?�U�hT�_���]w�3�J�䐔�4fW�d���������p��"��&�e#[dqzz/ (�\�{���S�I���N�ݭ}�уi���)�?�����z�G�Vػ�<�.̘�.��	7u�%r�͆nXQ���!ӣ>��5m��z��P�i����r��������Io��ph�әq��4+�> �f(}܁sY�ד��~�ZM����h]E��	��4�)o:�	��`�����3�=�#�нf��'�Ɔ#��	��T�:��+/p7[����n�	��,�>`?
�l��&�	$}���R'�j��q}�\�_rezAax܋����cq;�*\Vf�"/�eX5�1?\(�� ���Ԣ��{vJ݃Ss6/�Iŋ7��>5�J uBʺ�-[�x�\���b����g�_M��m�{�'����T�4�S�$��5�6j�����Fؾp7ǥP�� �*�?�s�L��
n��ZLH�^1��)ݬ���(�]+A����j�-t���ڳh�N9�`�93!��N����ѹ�^8�g WKhwɾ\��1�Y�������2ܧP�
瓛ބY��R�n,��<� ����'�P�Uޏnr/P�$��Y�ߊ�xû���k};B��D!�Ÿi��I��Q�1�^P|Zn�ī�o;B��e��fcM�e����Z̕��J�qz��
MrƤ�����M�z���ۯ�L����cn��e��mBZ���� ���Vk�f�k%�й���)aU���x�|E<��A�A�����_Ձ��B��l�yA��3r`=c#5�V�D�pǀ��ӰH��7����niu����K'^��w٦��m�H;c�`��'6,:�h�����T���ɕ�p�)}��Wĩ�.)��!rxu�U���9����/M�y�b���10���.
�=�]�(�&�9h��k��w���#�pkcs� z��(J����m��,���Ձ�S�6`W(�Oo+�Ff�����&�[^H�6�c�/X��%�w�*�,��Bh`@J��ž�v!B�N3��Y��E�!qF���3T���p8l�S��:C�4!p }ЅXwb*!�f+n!��~���x�^+��H�l�����T��̵*��4�d-����>b���QEq�����r�m~�2e$K[�3���ܤ ��ӣ,���ӧE*�i�Ӭ��x��¬�U�Uq�OR�_��Ⱥ�8��g�����P{��v=��{uhjpl+j��q��V�S�_�+y�|�_/=�g|������#<R%��j+�R{u�����H�to�C�)��J��5	�Pd1Z����:��9Զ%����:v���E랹�i�h@��߂�l�r��PE�� J��]�)qE����j�p�%�Ӈ��5,j�&qq�Zy���O�'7�W�z�xnt��ǁ��И���� 9���BO)����@����;�m�M�������h�dq�>M�Y?m�����O4���w���+����]�.#����p�.g3��2[j��أ:�%�a������t��Av�lԎ���bGºd7&�O��V�5�	j_����?炭�H�яs��H"�$Ŵ<���k���-����/X�w�*j�Q���j�a��UT�����^3�Ź�{$���5KV�`.*k�]d�($!�@'����+�d���Qj���B&O��Y�ɉּ�)��R1YS���=�ƒE�NK@�%!���"�c6P��5ԭ��K+&DW�h@�����v>2����� �*�_�LO��z���M��%�,uEM�ƫ�q;���*+��$�b8�o��=����KA�n���8�=J�L&)Yk��y��������>Gx�B��3A(7Q�ܨD>������:��?��ܿ �6x"�n���<t�#��W�����i�c�~�?!;nm�B\GJ��HЩdj���GR��,�
16���6��]�Oow ��ܵ�%�����]��Vм�t�"o�_��,��B��}H:`�yF���w���j�q�U�I|�����y���>��q$���DD�t��(a��vB�U��6N�ө7q�v.\W[�	cA<���7��Vʇ��v6�:��9�܀��Sx�"�[���;�.|0\��((��f�M���߃I�ryư:��.�I�a&��g��t��j>��vA���+t5"�]r̹/�B>ޝm<(��N�;Ű�G_��î=#��;0��TKd���p��V��hO`�	��<�h�Tπ6�j6�E�G5�mT�lo1�H�^�A��B����<t���8'�$�tŏ?3��n�8q�ȗ�H�S�r�
w��t��Py_��_1��OF'(��Ǥ������pQ�����5(�V�[v&��vi��c��0��q*�~썑�;�!�r�iҖMc0�w��Vh<k�2E\z]�`��:���!���2�q|C�nt����I��s��7�QO_�ۊ}�V�"k��S0�ݽc���Ӳ����f����oKc�
6��"�G/r:,���h�C����R���X	��O�B/�L��/������0lF�~��Z�0P݋e��Nk�`���O�ͯ�2�#�=����U�_�'ap�}	�`�/3�x�lZ~�Erw?>�������vP5K܂�B��h~h��%hJ���s���'�W5*�_�}�F��+�@�㻉�Df�m!��;��G�m�y��0������G�O�V:"��J+4-ȓKW1��Ǆ����!Nf/��%θ�����³Y�1�v�����`��A�ϩ���'d#��o����-��P�w���zGB(o��t�Ev\!W8/�0�H�O��{��	p�ҢI�����wTL��Xȃ)R�]���ꕕ��<XE�E�W���}�;�~������+a��9��s$�/�W�S��V����^��G���l���f_R@�[�jԈBNB��qP���*�]g ��Q�OQ�EC�X/�J�-�-P�U��E�
�4���j�@	�&������jNv�Vjߠc�O.���~q,�'���NWj�{���g�F A�Q�μbM����EO�l{���.�;]��{!Z�\�U�[&#���HcΔ/MyRb��{ ����;}g���y��K�Cu���n�ƈ��)%6M�:�ꓸ��#Qk��a�c������N���}��;5�U�ڀW@Y�%0����^��^�z���B��r�\ؠ��?@L��� ^R��d;�����/m�:�%�'�G���`F���a^<����?�?3{�uZ%t �~��xI����l���}$a���RY-��j��q �P��0��#NWGgy.Ȁ(����|��4 ��.���+6&��#n/��:����e)Ǯ΋T34! ��<ؼ��	ɮ+�g�0 �'S��Jiq�02�����*�Y7[�cyK�F7c�ΛS���#^|}i��3:&b�>����Y�ϧ
�|I�!r9wV�g֏ъ�]���Tȭ]e�ո: Sp�$+��O��AY���g�DN��f<�}��Xb����J��o��vE��@A�1:9�pp 5�9n�D;�&�����
������8�w�G����GbT��6�JPu*�%� y�f!K�5���}�u!a��ܟ̊�C�}�}�2�z��d��;*�yx)�frځy��+�͛e�0DF�v?��CFo����1yg*�c0��/ĕ�FՎ}��l�d���܌V�����a�*���vÇv�_v���&�6�� ��7�΀��3q��KG|-�K�K�ڏ��i��Yu"�t SĳuZ��6ܝ��}�ۧ���đߠW:�}8�柆?¿a�TA�a�1���~л�n�>�)���u���%�P��"���q�z]��	�x���A�x�Y,�:�X4�\q�3�%�|��ϛ�L��|������򧓁&4{�J�-R�^��sJ�v��Rq��Ð��W�;����⚮�a��[��s�oa�*N�q�>����wҳo�m�d�S�4�\7�ы�f�VUwt�4�������MhΈP�u�\�����|��iBݲ�δ���7�.����N����!���-ˡ�H�ct'�`�A�@��£z'�eȖ�'�x.[T-O���W.�]� |(�M������4�����
�x߰��f�7�Ŕ1���doq�Ȧ�~����?�ӽ5T��|p�@�F0	)��ګG�@FEL򛭋İ�l�*�����]����v}$
RMzJ�!��-���X��A�!��&�:d ��xs�Y�YH)����u��g��ߍ"6=Tހ� �!Z�t���c�P	t�UV)���ߡ����^pG�.��HQD���K>�|X`��h��7�X =S����
������R�w.��zNB�h+��S��l~L5W&ޘ|�9s��O��M����L,�M+�� �
o:c�B�yX�"�V<����W�Q/��GzNDe�^�;�{q�p7��eW�`!�j/�4a�4>.W�o�"�r��2������^���FN�n��X�D�x�T�u�ȍ�N��f� H)���`��}���d�d�4=�ڭ9R�3�P3X8�������v�J��a��z�/1�l[������A :IB��Z(R �1�c�_Q�2M�i��T���ط�����T��&��T8���T�se��ߑ��$9���ǎ+�~���pA9.
�f���I�{0[heD5B^J=�J����cZTg9<��<l��Z	��X|��JDt/����)4n ����qaEG�/w8H_����\��K���e+�dn�X¢�u�N��0
��І92ȅu�kS����U+#�Ԣ�>�Q�zѶo��z��+^�C����2�xx���v)���FWq0~uC}Wb�Qt�p/���-l�J���n�/��e!v �~R�i�d�x���o>(�x��\:��{Ⱦ͒gG���m��"v�������Ɗ]�ec[O�\�̐^sGQ���%�`����~�������� h��C>H1;���Z�>�=R�}$ו�+`�������o��a"����<��D����X��wD�'�B��W�d��㯐~C�_�r����"Tq�}�&OT-������	�h��}l��i���g�!�f�P�5�v�(�e���vn���B�KޕP;�QL�m�/%�3���(�����&4B�z>`����ؗ7��F�7��Q��be�@�W!=(���Yʱ�����$���|m�3/8�[�8�t�[����Dx��U-��� ��}��(��+��xZ�9�$�ta��-���+E�a P�m&T��ċ>���`Z4�i��K�U)��=ڈ�S��za����.�����U���T��5P����4��x����u���}hynkQT��sµ_��T��c�4�3M	Y��	�a#9���k�;H-��@�A�g��(���$��l�+º��h�A��E��5%�A�zL��o<K�C~������	�����M���*�*`Ӏqb.kw &P��-�#�y��s��T��{}���o�����㺏���<�a)K)j��C|��D�:���N ˂`���|b0��2�j-&��� a�_���Q�.��f4.N����h��B��St�T�n q�t<�5D�x��^�ҽh����&s�R���sނ�}���'�'k��а�;Q��JQT,.M��]�"����0��*��|�͊�^�� ֪>�/�8\�ʈ[���'���8$@);;ðj�,���RǱ������wU<���ndG�R qw}<wD>o���Ce��R��%fc�1}j��9ː��?0E1���
���>�5�V`}�]s,+�,a�c�]��0����?{I���K�B<�x�ȳ�I;���;��ؠxa�alh���Yu��#4�:f���U�f�J+��We��0 �G��Fhv$UVX��XB���>��V�����U���e$�:<J�q��y��G�t�W_%��q�(�Sy)���7Ҧ��E�%`6ޛ��Y�I��W\�5��\�0�J�7���lCu���Z�hG�.Y1-�H��̸�9 ��\�
�D��X��H�؟�}��9ś8�y��$Ȇ\O��34"�!��RW�e������"eY � �P��ǈ���-���K�+��o�;2Nu���16#VV+��4���A��*3��&��p�J� #��R���6�*�@�T����Gg�;�_,0�8�bϢ[����zZu�Q�A�1fHޛ�FWVZ*��4�R��3���/��<@�։c��#����$+�b��U����(�I|f*-���;˜[IK�*�s)�P���eQz,����i��N�^X�V�w���F�G�&��M�l.�*NBϲx�{�eĜ|*���:�eT�����P;�/�Ԉae�
���	�I�Kg�NR���S��^�3�ը?�K9�]$95����p�?;b�0�l��:��m���|j������	*��N���gj��`?�v�W�<�[|�p9��I� '!�w�����8���������m��N�p!��{����'�OPS���Z�l��]	��,���������̚�ff2�������'����\���&��e���X���l�&�h@8f�P���K+.w?'0h�v/0���M!��`���Y��G��!S����?IԼ�`���1~	Bmh	�65��8&��k��Qzk{����HnR�+K'��``ሾ>��P��ʉg�����,�ז�Es�뚪���5�*]�TD�h?�E��ԟie-����`�N+����T��p�F����'�s_�D9�z��)��Ĩ��e��n�` �,�\=�x��j�xX�m���8
�s9��BO��	���$yI�ט���d2
���&�z�f1�����W|4��SL8�K+�� %�j\a�n#`��;>#sE�=�Y5�ͭ!�}���jh��B�;!(R_m��~[q�6ƚ��Fn
�? �'kZu�g�9�c�Tw?L�T4��H>/��r#h���mG�n�|U�[�o>:�@m���+�k!Ph&e@�{�_Y����We��@�Lgߛk�+%�菹�p��vO�>8�:���mu-���u:��ɡϰ�p�ej�qy��l����$�Uf����_b�W;��l�M����CE`��-]�F�U�QD0��?j~p�W��5I���ae��9��fM�tf�܎j1����%y	��j:k'/Ϧ��KB�a�i��X����
*��X)A�$��nj�C\�$Y2i<S3�h�K/�Y1^&q���83r�B�	�
���~�j���Da��@ߏ5G��M�yՄ���{j&���>j1�]�ؑC/�Յ�1v�¬�N���Iگ|f��#��L��Z�S�P����tj`��vd^a� j��h#X#`�,�)��gMf�u�ZF��\��E^�p���sOyp/�Le:�#'ͅ����
�I�����x��@�f*"*�'T���E�(m�7ߍ��Ǔ���bdc�gL/y"J�\'��k�a8N��Rj�IKލ�p|=.�/y$c�d8��s�v!���m)XN9����ih���t8��E�����9���h�}`vo�9�R������W~(���']��q|��S�g?n��[�#SK�Y�Z���$m\ɳwu���5�����RB[x4(�7D�Ļ�5��gV�ew����TQ���Ԗ�k)ɥw�WT;�1e�hk�U挱!�ܡ��D�-��6��Zr{%���Q�s����� O��?���c�_��n��X��|�-q/�a�p�&#�];�pB�
(���_fx6ւ[�)M ��yWh+�(!A�p�:��d�o�t�<���[byB���P�+zQ��ׅ\;�f�<�Pm�:��x#"���/��*�,)��mh���}��������0�ڞ)/�T�U^����!b,�LIA����u�6|?�0^B.�\P�����1��-UbN�5�,8�����tR
o��:�DJ���� ��WĶ�}b��wh6�I
D�7
ю�n�)����籦���*��+�j��
c̜������e���G�܋tE���7]����*w���|��Џ����,1�Ϯ�U%�in��e2���>��*(�{��n���k�E�`qk�m���V�0=�1��q�*G��8cG�ћ��abm'R̂G�Ȋ��rD< �W�l��n���mӂ���2�q9�G�H�
��y���0K1sT��Oy~.`p��nw�M�ۙ5�A�{$(��� �kǖ�N���CǦ�<�k�e�@�9Q��2�t�y��SJ}��9|�h @QsƁB�ș�
���	~�A㏰����P�������G:�/��22
�
"T0��/�����9 ;k$V�ĉ�� �uB����*�,H��/���g��;�~�~�B,��$���a�ς�5 d�=�p�Y��U�GM y�2��^tʕ�=�2�J��o��Ʃ�C�k���.;�ƀv�y
v�i�?Y�tM�㕘E}`#�3��c<�#�seAE&\Q`�x��XO�a �&�-(k QW�v��k��I�w�4��	䓾��l�ү��8+���@������^.�֔��d�g}{󜘷��9��\�Ae����mW���F��f=d�����}�}'�Ĥ��N�@A��<$��m|a.��`��@�r������7W�X��UXԇ���G��\��Sm��T��c����`�Ԕʅ��G1Ϊ���A���eVsw���N�H���{eN������uMK�1� ��\_�W�����bN�^[���5(�'��&�*eĵ���,7=��L�����0�������n�N����9KZHi�D�sgy3s� *���<� B�A���lږ�aS��6J� ����烔g�W����3H)h�p#�Ր��xU�C(�@�M��P�t��%T����y���f�g�	Ĺ�_�Mc���^�#�x/U�7-���OA�ތ������}s�Mf�%.���+F�V.��c{nȸPD-nk{�[�w���>�
�"D����3c9�ʨ�:�Π١x�d\T'_FV�7偺�����aNx��	{���	�"�j�&�'�F���"�I*��,���<�w��
��V���){N,P� �H��L�j��c,h{��v-\���R$�	tK��D���[��<���e ӈR~j�X^u�.ԙDwn�����A0?�'�A5ԉ�+��x��	fb�nhX�2c�&u�'a��Qw� xX����`��EjW,��5�`�hl�ՙl���sw��^M�~����?5���S������Z����u;;/�A��^@��D�����7��XPW����_���7�*Ky�?���95HHN�=Њ�M���EN��"wJɭ�l������AG��)�ژSI_��'+�7I|y����D���Ď��Gh���ڽ�|�F��u>fPg�.9.Y�e��Q�4y�Of��H"�ǻEF����]�4J�lƃ��X*SP֦����?�%����hw�<A$V-QӔo�db q�
C�g���,7\�����!< �`XO��I+>�>�O�L���#��ɷ��O	�4؍����E� 0B&�t7�p�${���lk��n���Ak$A��z&��~�x��Ygo�ۖ_���\��"(L�(��b%��s�I��A�]���e��bwRD'�I�vw�D��(��b�'������r%xŀ^��j��G-�3�|�n�� D&6���Y��E%B�rF��`��S��mO
�M)[�ڱ���uc����`�ڐ��z#%�p�?�g���`oc�ӖkC���a\��*l�[B���Т��H^p/�̪S�h䍱iD�ö���*��5��Q�f�Ҩ*�1oRo�Aq3��$@�8���
���(�"�����_$|VQ�<�A"7	=<�H��Z:�]Sv���ޠb?>�Ҁ� �O,�JL=�����@��| `��S<b�1�)�a��u�N�i1�X���A�ѩ&�����{�Ն����0��A��R�OW�Y/p�3�n�P����`�"_��;=s�p�ч��o�A�lt���d��`�ai��qDY�L��;�J-f�-7������˄�I��K䣃U��E�W�և|�<.!�(7�{|<��+ mܘA�ʡCh~��k���v�N� ދ���	ѻ�d��i���E֪�ΊM�Ь7�TL:4,<Z�ȿ:���C�mӈ��ƛu�e_�w+g
+!�,��S�?�b������C3Eq��A�V�{d(]C����_[�Q���t����"��Qs��p\���η���ӄ/� �`�3�V���v_z\u2$�M���3��9��@׃�O��kC��c��H��ּ$�f�!~4�?����<X򣈃�)���v�$_���û�	g��R�G�o)[4�Ea�eƄ��^mt�:�hP}�`Dx�8��

EۮԬd�y�t��̊J���[\��<v�k&*�%͐��c���7fQdZ�9�c��c)7YN$�ma^��pE;h,M�?��E�o�3V�yu�I�(C���Z$2�[ Fq����I�{2H`�?$r%��[��<�����'ҝ.d��+Q7�V�Lqm���8a�RR�����8���c���7`4"�C{lĞ�"�[|#��P޻�b�G����6�l7t[Ļ�+V/�b$�i��A�TF5"�x��L��G[��@�����\LD�u/9,��r��L4pgȅ���C,�ڰқ[R;�f ���ys�\E��'��C�8v��NHL	Hьс��f�9�;+{�e>�
����|D����1V�g�\���0	Kp�x�J�M���^�a+~O�yIN���� ��ı�����$]�������S�JZfa����٬+�(�����~�|���E�`�ܻ9��(-��ő,Y�h`�[�����݆~M'�(y�m��;*�V��m3�ub��a����~��ޅ{~S�:[柌��,L��}A}s���-clU��j��xCML6u���ְ>T�B�2�'��yA�V�#��'��hȘ��(b��>�V�ܒdG�3���WӴ�'yc�wg�Y�YRn��52��mX�N�Y�/Tp���D^��\V^�}X�!Vܱ��A�A�GP����.��8����P��0���l�[��#�ځs>�6�oxJ���LSuH��
:��*b��IѲ�Jt�j��KdŜ޾���rbG�}�wq�j�5E�C�6��k�5�T7�x���t�3���sǟ�S��[{d�m�oj��z!��b�{6��8����F^���gN�ʓ���{EQU��Xv� KQ�IV)h��݃�����z�=n�w�X���,9����i�zq��f��+~c�8����i�4^R5vj�E#�P�˟��V�S�Au�p��)+�DPH.Z�h۹0(�%N�zع����*!�Y��}h�v���`[�H��N#-�<a
f�G����]�|�u�;�k���<
4p��v�/	4[�˭y�kې�y��Vmf���!�?�X���
�@J7�J ��_rW�Z��#���7�˃��-� �%�|����x�ҁ)�%��w���_',S}��<�4�L�q����ƪc�,�ᗧ��V|Fx���g�]�C���S5l��-+t��������A����5Զ}76�F���{Ro�oQA
vzj�̤�W|Õ��al��5AQupAB�g�l?YfxH,��J����p���`ƶV;�Ȕ�0f`�!�g%%0�X��{l�K��^M�y�s��B�_�X�o	k�,�����Q ���*�W�@t�=,���Y�����[�?�0NGG�f�fl��=hټ�̡�G�A�w�2�
����*�c���~�	�8wI*�&�	�ԋ�&[[]p���`��==W-��T�yԝ:+��ްy��X.���p�$�2Aiθ^ޣE��
����z�Cj�a;k3��?��#��qB����e6=��
Ꮲ�6�|9?
�И��M�5OhB�=ԑ��lq��y�b�[����z�V��s�D-QF�$��W.?���S��#�>����@�u̳< TO=��:%Kb����`� arp.H X�z�V�z��V����!):�-�I�ԃA����1���U�O�g�(��f��	�3T�Ò"уxM@��}MJ$i��H�i ��s�v��N*�ݷ��!�B��Cg�V�R �/�������@7mg�G���^�W�Tj#(E�	�+G�Y�)�5��<�e�#q�E.��T~7k���1��S	_��&C
]2q�ԑ�o�ޭJy�0��^�L�Y'a�����3��-=]L��S�M�������w�R�aD̉%GV3��=׾�m��s'�/���2lj[[���<i2椻ѨJE�K�����x�i���G�IAR(��:�ir�����Q��J:D�ɉ�@γ:�f:���B��N�]$b*\,�M�T�4��"#қ�b_�>���-�̈��i ܅�v��j;^~%��EJ0���D"ƗS�Vwx��L�?:�S!`��U���Ք"2=u��o����:�T.1��r�><�w`}(SG��ZQl��-4���&^���d���i��R甪uҟ�)f��,��E�0Mʗl%3C(j<NY��CH�X�Q��
�F����Ka-G'��/��},$������J�m1��P;L�^�I����K=n��KM�����Y��Bψk|�P�úUhK@���L=�H,S oAϬcf��̉��!i��cP�;����a�.kr��<P�Gr�f����h��r��B�`>֡���5�Il�|T�zӶi�;�������f~�����@��_�X�TˑI���4[��W�뾓���HXc��ǹn*g<q<���D�K�ջ6��M��|�����V��n������ ~KH*��&|�I�-�=*�|�o���PBG�C�e�c��c�/�$��%�`k{AqK��Ջ�kE{�Xo�]Ƀ�%�{��)������e�LJk]��a����H �\nq�m��m[8	B*��ۯC��7|K`I�ՙz��I�p�u�o�L���P�_?� ����0�s1��յ�J��9k-_	2J�ȴ��ĸ������͚c3�F�b�n˿ɰp�yF��;$)���AzsF,�I���8��ԅ[�?�Ϥ�fE�����&un$*f��i"r��4?�����r&���/��aHk.rl�ӝ�N�A��22����� �!���\	�}=�h�
��5��P�=!}�΋Jxw�t��[Gƫ�Oe��j�;B�Eo�Tdf��t�j�� 6j��C�)Ye����KS�+H���-�W�tܩ�V�nR�L߉H\�	歭����O��j
8�J��Y��N��VSw3���_:N	�Q�9�^Iq9���	[�>��T�i���њ�|p�Ē�'�����Ÿ�qfҘP�6�Ƨ6,n���w"=��K�(�V��/1��`6]p��Dt�D#_wPk�ц��^	}�嬐uG��쯖]��%KdJj�Z^]��Ӫ�~��bߑ��~����{��7~RǮ��`CP����VC6�s\��vQ4�AF�&$=�%n2�b�# �jA��=��Cf.�<��7Y���!!F�8 ��~�n�����TlO&e��bGڮ��ijПK9��`/iY��Ho�V�PD�Тo黻�=<�_�`#8w�
���%�ALy꒩������n��bt�YXBpV��i���([@��O�����K]�}��Å��ߩ��4�w�_c�^4�+��P����_=��g��<<��P��_��u^��I'Y��62�ZX�yD���V>�ev��.u�����b����Qa�o+��A<��?'����l{�t$(���*��d�J�_��:�F��6���Ց��D��Xi��}�g>��w����]t<�lB���#�l����2�1��ۥ���u���W� +�A�N^By���K;['t~��{%�����2�������Ȗ��[6d���k��c�d''�i�<�~��c���#�����6�+��ȫc�.��M�@��W�*:���s��u@��>�x�>h����k��Mn��U��^.֭�Ns����=#9<��L,�O��!x�`6��ޖ��q�ʼ�@�D��ҏ#v�{�z
G�	�2vrBJ�j��ָ�9�ţh7#WB�HB���5|,5X%	D��	$���4�r�Ծ)��/�ip�/��c��2}�K��iv(��bT�`�Y��Z΅Z�s��Pb�x���:\GX+�:��xx�V����� �:�������n�Î�!s���al�U�"������D��F�����[�1��E�>�����Qk�hʬ��;�p�R^����y��c?�0��;���mᜐ���R�z����;��=���1��������T+���a�|�������<����*����?+��՝ьK�&�}\�X�.�`���hK��'�՘q/�I�z���t�3�u<"���p�����u���@������\�<QP���P�\�y��JU�#�� �<T�
�Zk?&-�~�+�L�ə����F��ʱ�^��/��E���]�6�o��@$�'5�뜠g{��0b�-
�v/e
D�&ӛ
(:]\0�V�6bOՁ��	��	�o*��/� �|���urJhn��qɣ�+	��)�k
:�zK[5m��
���֏��3@�N�mV�s)���]�xq^zn�K�W5t�{#�t]��nL<�����Xg�՝ҭ��Zq;����IA�V�8f�W5���V~��t��q
/����G9�.���
��Pa�G��X@�� ;[fL��DQ��QȊ�W@�N�]��e�����*��IS
�J��P�1ʈ\�|��"������jm3�Od�i@R�e��Mծ��wvBdn�2E���[�/"��d���G7n�6m,�5wc��"k �u�8���v�{:�5�=�	���_7�C�M�:sV"�RW�
����
�ў��V�U��
�f��]��F��S��Ԓ��n�V�;�5�9�r�
d�����i�[�X���i��r��iRɃc�;�D�C�?���RA-
ƃ�K��j���_ȍ������Ҫ� ����c.�u�pe��n��FP���)إH���.����q���<C(�>B�;ڿ��N#��d��)�^������Q/�=zܫL�Ol**H��1W:�K�*��%���c*���b��=:a�M7��R �ƑIBf(�]݉����3[���A��u,�yfZ�s����< ��䲫��8��m_H(���9yB�fJ��ʗ>���'�Q��ݝ	���X��_�$�J1�1�� ��>?��M��^���=��k���A{�A�yޅj�Y���Eo����q�싉�0Iȉ�K�dJ�h"��u�we�c2����R焀� ��/n���uts8��H�n] Q֠+�(��y`kFl1bN����qڡ����8J��H�u�Ћ�[���nF*!�U3�H�?]��·쪢��5�3�S�"��L|燾YYoS���2_���h!�6te��h�w[A��4)e9[P�+�o�q�:��jq;Qe�Mi��m:m���r-�v!9$��=`hM$�Ɲ<�D@,*h����$��.��[�R`�9M�{���P��\~�SBp�*[�0{3���\�w��hr;_^`3G$�CL~�L�X�+���D�5-{�PE���C��|��_@~ro�Y ���Fİ;qi�Rm"�+UQ�����I���mH9��y�Pw8��Ku"��c�H,���*W���P�O�7)� �J����CFe�A���4��'n�̓���2���2�8��k�6<u���c�P�<l�?��9iM��%KS��)�"�j����ݭpgN���M�ڷ@���)�#��T�7�Q9�ڰ��W:j�l H�V���D|�n=��S�>�����4m��Qxa0R4N���뛗1=�&.B7��Q�����\�U���Ve�%1��Δ�������1E������k_0���h�:�*�~2��Х��+���+0�k��W�؉['�"�n������mz +zJ���5xy	
πR�JS�슖R�{ɻ�as�Q1�A��li]�Ǧ���:(��G/��[oՍ3*��c�TGB�;=��{����'��rP�������U�'����_c��Ğl��F��>�PJoȑS�vۧ�LL�!PWTtʒ=VB2�+,w!������{Zh�{�$	�C�|5�8o���&��X�ͫv¹Y�*�o	�>��~�ԣ���""F�?�����F�:(T[-:�lQ���[���Z�h���H��ϕq�?�?Km�}�2lX^cM��_�@���3����v��9�tw�k�"-]�:��AO'�%����hM�ln=�+ü��NV*���0�����w
3�O�!c-��&��Ǖ��{#BJ�#&r�¿�}��!�����z�L1�eg����~���pJ!U�K]�Dr���@wcL-d�m��9沰��� Z���'�̀��zG��l�;	:�&N�4�L;n�/ώԕB|[��,�7�DQx�L��7vQ.������B_y�M�q\�����8I��I+��.4�7~\��V��O��I:�Pe�ڟ|�AI��ÉR�rw_��Vw��n,�`/��uBѨ_��ԕ��]W�����i�w��g�8Lb�2A��O�Rl��]'�x\Y9�H���Iwxڏ���g���q�Aj��oI�Ad�wS�x�n~\���� ��l Wi�~��c�W�6dS���#��	Wr��gw��gr��l��[D�����JQ����5��]s9��R����tJF��`�3O�;X����{8)�xP�}Es�������~V�>.NJ3w=Cj�0-�����B��?XTi1�`9�<���a�����}'�7�R�(����ЀW��V� �_���*�y�X����ܺ�nU��V'�b�E�.4�3��6�!}s���6(Ts���*8]�v�e����v0x�S��D�ŉx5th|�q��`;��^lY�u��A2$\��N�]��������4As����r�D9� t5�q�ڕs���=^e'�u3ٚ�ܬ+T��OR��		;�����k��,�X�mW�"������1�}Hh��Մ@S�m6j]vM��CNm�ڷI�s&엨��C$G��yI>�;ƶɯqux5��miQn��Od_���QP�Ա#����U� +o�k݂�|h�@�8>���i����Ce�Z;�d�(>&����oO�Ѯ<U�?vx%�����/��^k��o�w�ڍ�k��7ٔ���c��_+JLqR�Y�� ���ْE�+/�wz�:~��o��
7�IY�đ �!�+�I��X3�j��upbv��	uJeFnS5���-S}�?X2�#�#:#�˴����P�3}�Ī;C��	@Al��m Z��E�^��3� ��� �,�k�>_VD������fɇ(��{�S�����#uQ��pQ!����Ԟ4Y���7iɋ:ʑl*��'� /$/�S7�Q?^U�m�i�2�w3Q��8�Ę��FQ9���ZMkQ�ޱ�A�~��g������D��:{uv�R�Y��=gF�ne�QӼ�3dY��$guL����E��&��"���vm�Cq�շp�]9y2��:����T��9@�4_RZ�2�(Y�)�%+2,��o�Ӓ�=��?QD�����4_ȧY�oS������ͽ^݃��R�8.��֕�&��B>qɇK������ �b��f�o�3o��k�ZĀD���ɥPl��@Ϋi/�l��]79'@Mᷔ	Kι���3�9g|��;U�H�7��s����W����EA���}�/�&��a����#��Ԧ��]�w=���Ɲ���)�U����|\f���<�qL��Hf��$R=1�����.>� A�n�es��<��6
V�CT�� ���<��4�@g�	��@_��l�]�7*�'K��M]�}c�3�?t��޾۬/�Jb֠���>v�E�����ɠe2<9�y�A��9ĢOB>�r��D�͋�eQ����Q��4;���|�;��RA�R���?�~�����s6u��h��h�![]u���4z6�Y5~b� �3n��K����J��N�b�����1����Ec{Eᡋ���'u�&�`B��R&�1{��+�=��;�����k�'`�����!���K>~
vU%���YbB��mh���>.�|Z.x	ؘ���5,P�d,l�88Y�$�5�X���V��MyG��LA4�fN<�$��;#cQ��g��~�%5;�:�d�@#q��f���h�����C�0�	����?�=�3�̾��9����<��t9+�r!^q��QjY�?���0��M�] ��������M�ב��N���ޡ�&�j��}�E!0#jў�]#Ɏ}5�kѦ ��e�m>s?*/���&�������q�;S�=�Q�0���/��'�%G`2W~֌�?�1�h���H,�5*��>�_�zq��*��o���ͯ|UI�V��\.�y�	q_��Zf�-��1=��˙��/h��"e���q]���]\�OyP1�=m#�cA�Z+K4�Ȑ��|�】~�^����r��#�t�#���jW�c]Cw�fوZ�����&��3%H3,��^����y8B�x攜����"J?c>3j��7C�ZJ��d�JY��Z_>i=�	J��:�BZ1��Pl�m�`ko�6��`tj���@�o�Z�L��5�-'.��ѡ�Rm�S
G�et��C���������3Q9.���D{B.�&�(��+TD�rЁ��]�.�p���t�-���:�5_\#m������Ħp9f�$��_��焎J��X�3�~�5������kk�g7��0��q]&<.#`p�N�\��`n��6|�Κx�+z^��Y�k��
̓��J�QQ�H���1,q�Tod��>A[�V�ȸ�X)m��6�L��D��ռ�5�l�H�a��B'��R/e[e�h0�E[��u8ԁ�~ϵ����ҥ�/����A}�ɼ�+��t��wD�33��FN�g`o��h�kMW��'�[�֜��j*��P%��q;�a�Y�3ߺ]d��Qoa�T|ŵ9��ՙ1Ǔ+�)��?���X�xy�0P��k��\�n�	�!C'�J��H��6m���	�}�FU�
󭉓�x�Pw��K�,�wy۞3�,�ܶ!����[�N0���~�O��ｂr\n�oWެ�M�����6ڤ�u�Bk��}kKJ�j9fPS�<���1N��GuBA�����|������t}]X.g�W3+��fS���q~� �iAƂ��/ݖ��$,��~U����I�I�oM�(
�����Z.����o0�Ɲ�8�P�oi�f 25��p����B�.��J�/pVoؽ�Tt�jP��r'���[M����?�%v��)��C������A��0�ާ�Vu��T�-��;��
n�p�2k(�uR7��t�i�κ��}��B��A�2�ؽ՟u�{A$)*y�#�}:L'���@���AP-��x��N,�:�� �ܗ���l@l����sql��O}\&���:�����v
�-,!۟�+W���njE=�T����@N�k���`B�R�gw�.ٳ��ۧ	`�����,�_ò�?,mU����b��l������̌��qes�.yw�N�@Z�5���e�D�PNs����)HZL(��ז[�3K�h�9��?Zp��-T���2Au'����Y�����ϴ��G�Wɾ�P)Mԣ"8������;�ie�fp+������5O��Mwsx���AQ��������t?T�Ȗ��X�3�G�����pK�3�.�IhrJGn�$!�g�+R&#�#�Ŝ�ku��,�}D�j7@�E�܏,?" "�>*�y5��<���!_<�p���׿�-W�w���]�	`�D�Е�Gx�sw�%̩d)4
G�$d���X�{9��f<���7��lV����w��H|p�6�E:{��M�����<�/%�߬�P~�LդN^��K���i����1�T�!��4l����o�j�rb��=����?zR]��� ��;[����f���i���E��[��{�"'r��?�2R$�%�H#-�L��Y��h���8�����T��m��Dw�2�K�+��ɬ�����58�����n�/׻���
�����%��p�`��o��3ng�9��C5��=�W���H�Cq\s��
N�$5"!����
p[�L�|�(��#e����M��K
�#�WVw!�#!pH��2C��h�Ü�^7��熵�n�c7��;��dK+���YqM�5(�L�+ە-�s�˧]f�{��Sy]��a��r�ح�>��x��ju�K���l��:�xG���%'}�W�lla��f�<f�m!4��ݜ��g��,-E� Jˑ���,�h��i�˻q� it�#��h�Oi.q`�F�E�N�d߸�y��0T��pbA�c܄s�ǰt22���~<\6>BاT���3�������H������L_�ZX;?���N�<n�Ah��9_0!)�0�.P����D{�(y� /�ձ�^� X�Ke����NN}�>0��oRv3��P�gPHQ��h���_v�kd����o6^�P����]����KWs$����/��`��WL5!�,���B�ŀ�0�NU�:�k��~�L[�s��g6V��w�V�m�����;t(���b�y2"�~��7 iV)U���R�9wTq4#����\�J��]��$p�&�`Yi8H�\��>�K���o��5�䥌SL��\�?�I�Y4W��@�����g��*%I�[��!~�e��ڇ܂w Ԉ&�M�H6�o�?Z� @�*�I�z��S���y��~��i_<�ms�iy��V�x�@�++���`�Q�)�D�j��\���<�v&�Z�ctO���|�}�8�(" ���B+�fR���D�T��_t9�۾1|t�q
ii�ᄯ�c��k"� �VW�Ƿ�_�لӔ�F{1�&SY%<�k��`?�9vUH��m�z��pWl�T;C,N �����3�O����  V}"2nP�>�P��i��V�����7ν[�qp 6X��M-��~eEw�N�=�qɀml8�7���O֍��j@*������ŷ�
�	�ҼH�x}�����smDS��3�>����z�3���c���hha���@�1���
f�� �yC�kB��J_l��vc��8;[��QJ��u��Mf,��6�2�����V�ˏ��)A��/[O&Ais�C��j��w�r��U?�� �-�������tO��w�2+!��-��O�1,��3���ē��p��ǭz��Q\��A��b��A k?�}��]#�@���u���:�}<,]��z�Q,��/���/��b���<����}l�C�:kX��Ws�l�5���zXF��eY�<LK�EqE>��ʷw;�Z��cٹ��w}::+jx��Cqu|�
���Pc���k��zZ�ZtDX�9q�׍bhk�H�gp��U�ըZG���	������x�d�.Rm
N-�B�RB����ppk��(�����tez{�z��j����u�ɕ?$(����	��AZ_!K3�����w� Qn�~�v� �������U+m)}$�F�#Hؠ�m��b�1���ͻ\�b��L(<��<w)p���l�d���u{�tK]0��B�7x&��D��+[��_���F	'U�r�	��3�b&��I�v��C�j��o)ש=����[�RV��=��-̪%���4�p�P�A��h&�75�x&z�|3E
���֎�dG3��8Ԓ_�H���ì��b�f���K'�����q=M}%6�{c��H3aE���}I�V�_��l��W7��ױ}�]����;��Zқ��T��T�$c���z�M� ��.xD&����5ԫa���HL�+�HA��/]&�4��mi628gb;+����2�_����F-��V�0�8�z�P�{삆��!��sw����	�I�e�c���!�Z�a���iE���B���	 �Q�yr�<O����3@�Ӗ*�WK��i/=+4�S���!�z|�V�NyT���p!kJ�I��}V@�T���G1�V)���i�i�����qO��lm�;�N�
�������zFA��*]�x ��8i)IT�C�"�D H,�٨CX����p3��x�(����3}��'�ae��'~/���Ǳ�y�C�Jl���aU	߷>�v0����-M���� �C��ߍ*2�ÜX�h"t?ؓ�. �u�zb�3Ť�����r��_���&��CuĘ�J��u-z�295���0H��
B^���&v���x�X����T�B�)S�-�N�tI�^�Wz�]*]����j�p�F#8K����9��Ɇ��$N�	����>PF���m������zY�/?��ĎAݐ*��2���>�z����$�Qʵ��N�r���3���%�^V��>��*C��̔�%���T7��;-B���;,7bdr~�kA�$�V'#*�J^��q��iZ��vcpx�c>A�[��N�p6 ]�-*#���ׂke+��HƲ`o�mc/�y��f�D��ۋB��"շ�n�X��_�dSv(z�j��ms+�����2	Iޮ���*����ӫ���{1s��E��C�v����gbw�z%? fKmK�������ە	�����f`W2����R�"p��O�1�;"�sZ�דz�¡�n�<�oJH�V7�/�Ƙ�x*���~�.�3�&�Ϲ�&w��	�?��}Lj��� 2�T7|��d��C�1��k�����-zgdo�7�G��RM��[�y	w1�,SJ²��sN�����jP�e���s��e<��q�HJ�� ��5���)�D�B�`ۓ�e���ZIt��k�5�ӄ�Ά_��j�>��y��7hRIs�!g��t��R���ճ؋��ydFl�����*	�����F�8\���B��;n��$��:��RR\��Q�È����ʱz�^Q���~��=�<����A�����)]�t7 "ߘW7xZC��s,*��s-~����fm��'�U�is�k�*���j�`I}&�ҩ�-һJ���鿲� >q���n1N�����TӂzH}#�N��iik�����M|w~R=��F�T�3��Q�0��t�P�f�
�uk�j�
˗�đ�8���H@7n>؇rT_��-��£@�C�ss�NQ)�?7��N��<p�9Ժ}��Eo��!�YXIV`��0�r�	�J;�0�̇�'ad$]ޮ(����P�>͘��b�:.HA��%�'�g���XZ�"��4a3����ʛy뮔���3Gi��'��Q
0=�N�S��*I-떲�#���Gˤװ�u������`,N9�AL�t�7%sݳ�	=^J+ҩ֚��ԧ=˶G�Z�+f�P$9�>��F1�[�Q���b���?����BZ!�H�@���tB�`?u��M� C���V�
������$9����p��fi��6B�jK�>|7
�LW�]�%�*qz�S�oj	TXE�ظV�m�=bh(�	��(�ĹݘA�׼�-.�]�ۇ�j�t�^.�J�ŰbWA�)�Q�AH��F��J�K�BvϹ�y"��(C�d�lA5��_e�{��yܡ��Ri��}B�]� z��<�W�{�O���1� �7�i�R��ͪ� gOm�R-�R�8��J&9���h�+������L�f�d���8s����1-3*��y;�ՠ��pI���&�8��*ČJ<Rg�*] !Ce��!�q�)������]�d�r�uL�1X�W0�cG(��f�-�Bp*6!���]��nw5Y]z�.�P�E{���X�m$��d��A���<�+0����8���O�ɳ�OL�i\��%�H�*�:�ᕺE-u�G`����OԼ���uo1l��������v���C|��{m���?> ��m�Kt�?u�����)�$��&�X��zZWil����S39��m�n�nL'_[���Jj�SF�W�D܃"�x�( �89����-��T^uÓ`���ˇ�y5���|�)Ug�����Y� �o,I<�Y�h�ԋ$x����#n�1%]���dv��9�A]�D��|_ۍ�3�(��렶�5G,tNWNBeJ��\��Bq�����ey; R�7 �R�S=�p�#�4�'ք���6ԙ>�Q��߱(!]�c�if+��Ԧ��A�����m�D0ߞ��r�=���4g��$�2M���+����gK��G�E��_]/J&��jGe�e�qH|�!�6�ڶ��]8��%_5j�ŗrFݣ��ݦ&oD���OG�*�d�/�v��r�`8|^�#���Щ��~{/��19p��)��H	�5�o����+���v,�U1}�q�]%	�ٕҼ�A�W��)c��;@�1�R�^��L}�nbDp�}��#I�TD���n3�=[u��#l�&=���S'��ZK6�4l�h���Nk0���|�E�#G<4h������"�.��<��U.9g5e��d��
��&n�K�ZZ%�3��|��i+P6�s�zc_+��tcf2���?[l�Ո�R��w��Ȫ�h�$F)�
+�N�������BM���)Lj��^G��J���\�+����*���c��w5q����iB�+1�b��V�8��d1�h��-�����[,p��7�ڈ�dN�wǦ��w#կR�Ҫ�܉�)
kos��yĕ�E��Fԅ�������r�x�[7�N���eȾ�<�U�%@r^&�]���t�%+�^�� �QT���o�f��G��J	K?��H*�hErD�Ĺ|֓�7��<b�|�{�x����'<Y+��!��|xv)�uE���@�V4��Wx���>F3+�	��yx���'2]�����˃l"t�H���N �a�#h��F�p��=��u���*Ͼ!��<y����6���h1�ү��X�J��*i7m�EP�8(r��}��\{�h���"��҉*��T}���{�\�~�.%��$�Fr=Ȍ��N��e�����0ht�IeП����+}��+�{�`U�8�����n�%��W���Ыz^���.N�O�W��8�,�s�����o	���-?��査R���?�Rq�uE�׉K�w2d�j��a�a�4h��0Y|�����T�^�N���mˊ�����"^��2��wS �
'W2ͳ�)�MI�r5B�|1�?�i�*V���'��\g����&���:Ҥ�{-��lc�����H��g�p�h7+/����o��Kq!-��BF1�E
��\&��u�Ƭ'������X}G�^�	�f1�� 1C�˼.8&�aO���;|߂3�z*K-����	e´-	�% SH��sR�ߠ��?8sd���ѓRA��p;�<���A����WPt��:�	E�縳�O˾�aPϹd�2�����)w4���*�����n��fdW_�������-o�'����q�@a��QI��F%�cP`���d𱿆�(��}ނX[5;�����¹�*R�V,����.��f�d3i_��<�HU��nv���tJT���o�ݾ�/��xt=�{�N'~���h=r<w�K4��>bF��~�+�B�$�W��f)�r��M�#�L���B���X�H���s�+2��fwg�n�68�sP8T�[��o��h�:��`�E��=���G�������0��B�r��ӎ������A��<d�9@�Le�"^��7���vȼ�����1��f�Y��P����tÙ:Vn�	9m�e�Ԯ�>��'�l�}�J��� �]��wF��N|,�ُCu��2��m�v���/W��k2�p�hkY�������]�I�M.;���Awh#a� $*�( �&��-u:�������OG�8_��}k{}'_�=�����������0�i��D+�.`��^ds�2B�:a�nHS.&2�%Us�aX�?��i#��ؔS0�O�:}��2/�Bz0��c���g�l�4�����-Jq7	Z�� �� =5/z1<<�Pl�w%��Ͽ#��ҘT[� '-�.��&���A8M\LlTeqi������eaZ��]��1(ݕ;F\���/�	K��~��'�i�5�E��|�qZ<M"O��]��N���ZL���tsI�K
�Aq����dn(?2�\2XF]�<�{��c[��V���J�2��VZ�\�\�+*2=���G�!���6\�����@��KWr�?l+k���^�R[7,7!�G9<S֍�ޛ��6��DO��v|��A4����D��-%�"΀Zt#�	��q����;ָBڽ�~H��ZYZ���.��_Z�H%~ /�I���F'<��Į���+Y�.E�B�la'��I���,5��\�A����Y	f����/�+ f-��5�`��>g!ϡ9��O�EbѴR���d�r���$��G;��.�m���yV���-��%^9��Ds"�����j�B̻�SO���L���]���r�vLOg�$���9� ��v��ϥvKu���6gӼŤG����v�����x��N��0���&�=�
ބ���i�r+�������Y}؃A���C!����)��.�Xl1ߔB��G�Z3�5~�p<(zk����{�K�E�@P�c�h`�U\(�5w����dYVE]�ý�Fٟ�Wv�ui�i�Ik�v�j5H::'�wk���ݟ���(�]��ؓ��
 4A�8� �C?��ڌ�r��8 ε���ר���=��7 ��{�`J>G�:�Y3�μ��S[���-�� �Ϊ�r=%E��9����@�����80Ӽ�)��Z�Έ��{�����v0֨6����:��d#�j��r�B�(�U%����P�h/��V�߾��4h׾U�B�s򻚯���v~�s.퐦����0���4�24�b�����%�p��rV*�ʇye�+��G�(!��K�U��N���M3FB�'��D�+q�&(e
��a�|#D��0׵��:��H6������W:�ys?�āQP�-��Ubhs�\OD�-�e:{���P��U����\�}yI�g��W��ʼVDE��X`��h(!~b=�V�����������&��:��⢯x���m�-au\���G��S̆x�����J|�|/D�+jho,��6_��v�O����4[8�y�����c�%�Q�=_m�+v�wHj�G���2�0n��@���M��ɿ�t�D��(�pa�$������>Ư��u���ʓ)�/w�V찓L7
^�d
r!�_��uUj��m�V��5U��4�Z��|Tf��-֭1 �����5���=z���>�ܲY���c�}��83ڰ�LN�B�4�N���H�%fM�v�3�%^�FV�����Cڭ�F��y���Ԅ�9H(Z��@y�;���'ks\���ޥNZ�m$9}qU3l�v�P&���'���U|I-5��"u��H��u)`�T���xa'B(T��;R��A���s���VD�"j2W��)��ߒ�A>1�e�t�����i�-��� 
�Q��>��:Y̎A�1w�b{����~㰅t֜�51й�%")����2�r���`�L{�>�Bq�ha����s��`�f���GE��;���N�o��q��o�SrS�5�d���-���&�x��m�3yT	��u�Uo�Q�v�RVo��K����:'�� �������5V"���m�4�W6�6���H��x�8��\;M�0����� � UMK�]�]��[��c�p	�uK{����R���PA���K$zy�rĴ5�{���� $0s�A��6Q�28_/u*���Vo���j���=/O�A����e����xl��� �fP&AS"�ȓlw���b�ӝ��9�g�c��j"�8����%�ELoeyN�&�<@l���p�Tۛ⧤FĔ㦣�k��Ø�K��f�oAx�K�ı�rMb
�lN���m�Úy���j����A�{O���FeT�t�L�i�9�5a#����R�t�!�iA�I��,RI�ɄQ��3�d�~��OB��P���.�}�ahGŅ"�\�v�

�l�ݣK���T����~prS��2�~���x�Y��w�M\�3ۭx	S�'$_8H����:�X':�̫�<�)�q����mL~�ə���̫BLF1��7Ʌݨd����(M6�-�H �:^�`=AM�d1��;W\�̮�;�����݋Gl���_��Z�`��ўR�sD��{:&���j_���4��4L�������4���҃闉���Y:�$�:�^�a9��{��I�ȖI~�3\����~тA�W�q�nn�~������� �l/���F�'�,�|I�)X>{�PE��md/�'}�qo�8��ѳ��Mm��]X�(�1��4�O�e]���KU��7�]��5I�WN<�5��	��\ �r#^�@ȏ�8��4N�y^�_:���fy�|.ҙi�!����\�Ճ��p5�}P�����T�.��Ћ���F���F��yY@!G���ݨ�r���⊣�Yc��~�FB�����x�q��]��U{��R��T�'#/M�Uh���r
�t�gb�Ms2���N�;Ovw�z�)��g��(�~�P<���md�9cؑNdQ���Aڳ�jѡ<�/~
�zNB�=���Y������ԗ�_"��]w@4������sd8Ȁ�8U1���S���� rdlg�'�&������z�&����c�S4 ��#Dk��g8}�b�ӏ;��Tv2�p��}����E8�2��H�{h;%�
Z�7��2Ѷ--����gt8�$T)W�cgHj�S
���伪�* O/i^"�E,R`��\��T��б��V�ySݢ�J��yG���l���[�>�_�Z^��m�keTk��(�ϔ	 ^��.`	�ȯ2�%�JTĞ������f����7�ҥM��U?)�#�����qx��H'�k��Mfs).^̓�E�ՠF���诟��eyx�[P�0>�æFd���|g/q�U���Hn�!�i����Ȩ���|@�{]�J�mJtb�����Iڈ��#=6�ӎ�rj�B����q�Y��s���8�]k�)� �6.Z��ܶ�Q�"�Ye}�mhyi� �!���x����
KX��ɥ`!r�A�TE�~�5n2�(ѕ2��@xͥ��>W�$��)ΞJ/�ؗ(�3����-��pL�_��jߝ7ĥ�bN�E[��|F`���w;���j}�.q��Jx���t<���&t`�n��uR}`Q߄�Z��y��n4�������R܍��$ēe��C��+�Wǂj�+72@��}��nm�*xĔ��&�9�Z����	��?bӏ������M���0�N�R��e�h�{;�Ի�$�J089�<j��p�����=0�~?)9 41rH�n ��>�&�|�$�T�O7���E����!f47���ג����w�gh4��s��<-j΄��)̐l�ZZ���C��I�`z�C����ގY���QN�i��_��#̄��\jǃ����
D�tmS�����P�*K˪J!��G�{ZE���z����c�n�n
�X�ѭ�;�	Y��pY+\5�h�0���H+��{B�9P�f+gm��{fC�v	�D�o�d����ؙ��E�i�� ��Ul.�����m�����	�CM#��u�U#>��0O�1��oXH��:��G���6��t�-�#,��~�?]랧7��a�b��6��/�C��0��I.�6�k��I���T�$���`tF���u���|�.N�t�@���S�<c#��U4"[JDO���V����h�/�H�?n��
�P�E�/e#�#N�RM���N���v��P�%��18�|�fb�{p��MG�<�f�qw�au0{�� ��[!�-U����}�|�&L�0�� ���_���W��\�?����l��.���h�q�$�d�Rw���|�F�*�%b�BiO]t�&����"4x�'w_B��\����r�!�69>���d��NԌ���潆Ŕ��w�}�Λv S9� ���|��ۈ<����*����@�F�r�O�0}�0��4���G@�����ٿu�W|��G��o$�+i��#H^܋���W�R���������bx!�˓\s_���->{t��I1g�^���>�_��=���X}1��N��#۵�pbC�.<�-���&��W^)h�Γ���)g\�;��eE�a��l���/&�ZE��+��[*,���ĩ���R�	��7$�7</����d�~z����14��騢?�h�G�݇m!�-�I-��t���@���Ғ7�&��*���,W�1� A��+�����1���T<�1�t�V�G�Tz4$"h��z�.+"�������O��������e9@�ZEL/4kW��'1�X#C�!���ؔ:.{�x^�2N�,6J]`6bB�l�9��1��S�f�&�g8'�����K�����M���ThI/~���J#����*�ą`f���%��#�T�<%��ұW� ���%rʂK٢����X��#H$גMX�~��0��� ���Q[ȩHy�p���B��]�Y�23!w� Y�Е����Z�^f�%�v膷]�V�D+��ss<�Lߜ�>M��B�1,��|��?�D��C�Uһ�ad�u�a���C�Y}���&��N����|a�?�������C"����4��_���ȋ�u��n�f���A���G�\a���1i8���)��,+�S�5d�͐��j���p㒃�2��� �b�,�� 7�<<���t:�ȧ>�%��	��C�㢛�����~4jC�e���k4�#���+�i�Ub�]�6Us&ِ��k6��t�$Զ�������1B5� L_"�m��D��5�ŏ���H!Ҥ#R��iM��@NYB��tSy ܽ�:"�\:X'���׍˦m�<�� q�"6�SC	�<nE�̋��Y�ϑ|�N��n3"� +���B��f��#�1xZ��}�y&����z��/��s�\!6���H�o=w�����/�k�Иz��u��,i�b G�~����v)��a���V}�����{Â�(���c��χ�V��{F ;������ �ڈE&�]1'8��ˡ5�sp��A�8����saA�-�B�����'���X�1&|��Q��zy���������iZ���V����'�����rg�vh۝ZʯɆ~}hO&�_L��3[0�~h��YX�� �W�i�p�3^p��~x�`���|E�Wת2I�r(�R��=jS��T���N�ce+O#�9I��䴎�(�$I}��w6�'�I4L$	\yo,f�t����H���NlY;����%�l�e�=J�$�Z4��?��:5<|6���t���hP$���ձC�/9�E�����Z����X:�6�yn��y�m�Rd5{?� ,�3H\qɜ�Y�+�j���:���!]����Ui�:#X#H!s�˽C��Y���i����ى)wBH/��*>h bX���w�5c��L�~pW������9�$K� b�� +T9��+i����TV#O���3�����zrw߶z�f�F~4��=F���4bzՔ�	A}�N�z{uc��ś��Ig'�G������0+Q43�J��T�P��L��� ��.=Q�oej ���
���׺�$Ew'ޯgR�. P�Aq�Zg���p��ROK��1�	1�l/�����.|K�|`�Z���ӆ�;�s�񅎝e�D%����L�>�c��K�\���tj�|��a�<!��TOU��mK�������0_Ζ�C��!��Y�3�t�2Z�j^��{�����݁a�J��}DS^/�z|��M����.��}t237^��}����jh��g���O�{�^!�ZN}�cV����.)C�t�.OCsf��j]~��]6�s��ri$�]E`R��:Y�h�H�h���)�W��fB�p�)�~z$����<�>O�<�й,`J��?<H#��F'NQ[�4�\&�?}/UN"#4����<���}i�&g�^��
����
�����bE���Ҷ�da�X��jƔwh�չ�i��4BOYA\fL�tt�Ug�@�{�`���N{�7�槺�f"�k���=}�s=��-��X�}�"u������҈[��� (u(�s/s�Vn�]���Hv��l\RY����Wc����`M@��+}^�ǘ
�)���$����~��9��-�/�L�Y���'�u/'i�b�Ј��K���0+ i�cc�q7b~�Y���i��� 4�5� Qf2M)��d�}��=t�E�8ɲG���Aj�w�� W/�_Q 0`/�@	���z��*��"���'SF��`ޭ2� H�,Bш���l9��n�NĒ��Lhk`��qR�$G���z4�|�]���42�+svw�F�W.q��z%/�|���sQG!�}��t�Շ�XV,�0 ?�{�H����V�­���xXl�5�&���s0mEڵD���!zS!��<ȮE�N�Yf4=9����*x`Ss�Гg��a->�''7%���I��vF��8��J�m�h4�K�D���,�$.[������7'�sө���"�e4Z\��M���΃�����k��� t�2󡷠Y ������LX	�Z����D={iX�7d.�+�ٸ�F)Z?�b����^�K%sҔ��S�����i ,L��c`#��J���-%n?��z��L;��a�<�:����8׻L�û�gI�dL��]�_��q���G%�.�ڻI���88�<����X8qT��g{90Sʀ�D�)k�ڻ�M.�	���4�>ؕ3M�j�d� _-p&K�Ƕ4�c�N��#5�Lml���_�'�0!x@s�sWrt�����UC�{��jF>${sL�{������V蘻+����HR_�_�d��"����B�E��C��/(�Ӵ��'�D��ڭl]ҷ�'y��16(��ә/�S�O%�N�f�i���KmieI�5��e�*7<�:d�>QM���Z��Sg�n䀮����M�[X��h�ڃ"9:�S����my9�Y�-j3�����t+Q��эq
6�K�-�9�$�����6��`-��4���9E���*<u�,-�T���O���7-չ�������)T�;׀�r)����
�6�a(�7� ��Y�>V�L����ߓ�I�d�l�%�8A��W��$����#��K��a��A �Ũ�r]�r�#��ZꏌT��c(�Fj�.�o\m�l���oh�<�m�i�Z�ҕ�AѬ���V�q�+mJ�B��էo��^�*�\2w5{����%�N�^�E������=�P,~����C1p���<��g)
#�աNj7�hZ��=��uϋS6�����8��U4����X3��6>=�����(8�j=y�ޘ��<�xE�s#d�1 �����lZ������E-M�i.�,n�2�a�&�����n���`Ɏ��N�=[��
Y*���	@DB�-pe.�)2�uOAԙ$c�ٯ�_��l�o"���.��7���=�W���x�h�4v�RBu|��p�`%G1��t�/�	���녨q'W��K����C� �Av(y[q"E�,�S�m=ѧ�nG�vWW�	sӾ�R�Q��C"�㮝==@.ݦ��A��됦R���*D+x��n��*g󱑂�lf���	��--�&�:(j仜���!f��zy\U�9#�uݼ�tq$dM�t���I<�z2���"��"� J]�8p�).���&�Hs���A�ע>�5i2 S._6���J$�E�!~���.hA�y�W)\Q�J��/��$<���v��nQNz�3[� Csv"|�
�9��1��e�~it�c��s�#+��Z(6��	�믵K?+�
���eq����4F�8m�����<ȇ��9��'X���b���q����O
yzHoQ��Z��&���������&���y'F��Ȓ�-8=�j!B�EA�r�,�+��E�'��n(ġ.�1Q�:[��>�"��Z�d��q>���t���\a�eâ�:q2�A���p޽T���]d(/ ��H�W�G2�ц������eZ�'�eֲa��=�����/<��?�>22i���L*���@�=Q�<g��z��_-��a���@3$~�*��b��	�Kğh-f�a��$�C5��HΨ������)e-�.%l��3����3�A�t�NJX+pK���g�f�[F��`��T�'�$5��r��O��γ=6V4�ۻ�GGJ�
	1��Ca�3 �t�r��gds�{.g����iFO��ɰ�Y�K�'*�$$� �#��"�P��=�DX�F2ɘOY��U���?Yr���H�-v��`�MB����d��fT�庇f�����y���_m��ø�?�Cs-��;Oam�AS�U�o�7�3�XK��7��>D0�}�NL9��X^��	��"m��ӑU�W��\"�I��K�dm�/��ي�:�Ry��ܤ5V�gt�Fs�b��?�ĕz��^~�V$ʂ�|���T���9B��#��A�R��E.������1!���XlI
��`a�i>@6U��NN�)��rd� $b���qq9X��ϵ�
K�ŵ����PK�*�J����=OE��.&4}���K��M���*���;����X���`�㯡��b�me2�.RT�h"�B�	��9}L��$���{%�X�V>3pħ�P�Zx��A�嘆��Js�j{1��}�A�1�T�,��/�i����9q����q��eE/�K�z�G�Q�Ȇj%��k�6z����?�?k�w�N�����cy"#AK����
���x5O�f��8ԩYS|���-����@�C-���R��%�4cY�t�4�����R.@,E��>�K�~�'^?�52Zn��7Q{�aD���>S�b� ����ȦgI���Ǐ�vON�I�T�#ӞVW6�)�rL�SEٛ� Lx@�r�n����	�(�Kٵj��?�S3�jg*F~�#tA���e�ʛO��=OzE}��ο==[�0�>�� �b��|��}1�/����<5�@�� �.��F�@�Ћ��xZN�D���e3.�x{�xC�QW%�l��G��Ϋ�d�g�6� fe<^`�����,��}��2}w���1�쒲Q�(��CE�~��ȏ��|C�~?$;d
R����:����g7ڪ�<b_pS%ֈ�^���[jہ���|N~%@�����x�t��J�YT=�T�����F��@��u��bhдH�����u;6�������Wc.)Z0� \���X��<���Ф���*
q.Uh�OuP����4���H˲ ,�������#`��v�Q��T4�����}q@�W�~�k�[ �#A,�}6�5S�׌/�Ʃ��||-#�Hz.N-���z�+7I��A�������ّ.�����:8����}��P���9��k_/P�"����m�p�n�� y���!�"���x�$��3�v��U�a0��� �w�(�/e��b��J���o��bXQ:6�T$t|��fq��`�e�G���3��O��1�>��_��p5��7�lYO�p"*�n5�ph<��������-��<��U��c}9c�= ������ĺ��0�K���9RUt=j�_�X� ����F@�a+�>��RKc�]��Qy����v���L�0��;��>V�X�Fy~l4���x��
�)� �l�-6�m���.�ڭ+�$4�Y��e���
��X��3���c�Z��?�ŏ˷
Fz��Tx�s�n�]��n�����6��dK�a?zz��ۨ�zSg�|->���ihB���`ʎ�2C�����7��<�@Ò!"��z�D���� K�Ũ��0'�\��&�����ŹT��bmytpףk?�lu�������r&��fsC�x\N{�V�ϖ�����0�!5 h�K�~I�RR3�S���t!mg�Y�>� p˻�O��%�N��Q8B���5��{������:ۺ7VD��E>�@"wg���ŗ2�bGa���\�8�.h�zI|��r�Wy�;_?�-��ل6���B4D%��[��D��)(�@�>=�ڸ���������������V6Ǡ����&�:���ހKjS�> l�F���"Z��'�	����[`MGDj�B���|�Ej<Y��AP'���RWa��%n�ϦҒQj�֕i�5�H�l?�v�]��]����h!��DT*�ڬU٘S�@�+�(���k+M�:7�԰�^' ��ӛE��~��|1�D��g�k̉xx-���|O��B���?�G�ݽ5d�l���� ��#¾��;p�.u�(��?� Z�d�U�k��T��J�L��l��P^�B�h�/K�Zu�h(�D��W���5#�����i�:�1|�Ѡ���.�a�������B^	�T�nB��:��,�<ؑ��x}��R.ϖ�wf>�nN�g+=���Z���@�[.�!���s=[���{`.��\z�IP�̒r���+HMzݵ
��p�.d����7�u�6��;���ܾҒ�W�(��u�/��u��E@��U�Ax�Ɯ�nh�^8�,��O�H	�(	�p��]��<b�4������Dcu�T����@ۙ�c_���������x�hJ�I��S/�r�r�Y9�P_c#�gRQ{#�Z^Kۢ�3Fw�5�;6;\��xƏ�M/xؒ�(BD'}ۈ�EKH�!?Y��9��#�xY�ާ�����4��A��Kzk�����ŋ�����P6�*!8&�r����%�`MW��y<�*`<lD)�:�7ejUK�w�:僣�m��fvP��z�]���񖌝g��U���T�m����o�q�Ρ>����}^u�C�9Y�E-=+���en� r�hʒ�$�[,˷�G��
{l����ϑ��ܺĉ]�$�7�T|�~UB3���b����GˉXe�֞WW6����p۰�)p�`5!�� �
�P�+��/���B��~�=����l�_-h�r fOFO9�4�`X�2!�E)�'I����X�^S�,ɷ0��Ω����"��i��Yo��PvF��5}b#dǩ��S�P-hA�a8�������(�{�rv�r��BJf��x3��B?M�eHEں �7ܚ\x����� �Lf�q$�p7��JQ�|�;'���⛗M(R]�����/;��I��%�����vv���fMvj�;l��h��c�����A^�O�6��0\Q�^<��[Lm&�����_@��(�}j�r�O���s��Ӓ;Lyu;
�_V-͎��1�鼤�����m	َ�w<������'�����Jn�t�t"�1��3-Z���yY���7@dp���U�^R�U�;�& �������B��S������p~��x�RRBJ=�1~X90r���J��ÖP��8��FM�E�-}�,����;
-����Ɛ߉)*�d$`������.y����e9�pWʫ7�k�2��$L�����O���f?�3��Ŗ^5x�"O��h�p�} �X�^�b���ژY��bp���/N�ʋeg���f������:@~?��H0Ie=:A ��i�?7{kp��FA�����2�"�H&�q
(�=�;(h�ۗ�e����m��A��&�U=vߊ�i�?�ͪ1J?�����+��ϧ!��+�D?�qN~'�S>���QT�4EYh��~�,�^�P�y7�u����)��.��@8���-g�7Og�7񜈬��d���dm���@�u ��c\4�N9��B��ҋ����ߖ -l�!P)���J6A�û$���!jl�AXQ�ߙ�,�����l`zR�a����4������Ǒ�XQg8�o����X�y�����ͦ�����U\N�Ni�奆i�7�|���`\-<�P����J����^°*y/Z�cR`��1�/O��E�l_��.eBN."���~�����n�m�ͪ7d��?�-6��n�K:�0�
���������l
b��M���V�(A/-ȵ|����J�lL�8�� �H�ZW��{�V���F����]0����\��'���#�[������jJ�a�F�����E��hu��IH�����)���t�G��9b�oO(k��2�N���F�}�(����z:PZ�S��k�%IWE˂������SX�Çn���Ac\���Ի�%�ڌ��y��;uJ�ܡG�.s�'���ګ��s��NY�r�����E��8��&�����JMQ� �WtxT�a-3�Z��W�-%��<ޱ�'̃�A�+G�������wB�����-w2��spCw�EK <�U��(�W�Zn,A�6�Pz^k������(�"�J���!�"���V�۹�U}0�qe"m���=�"[r�`O����6�1�S�� o��o�ë���)֯�A��};�z:���i��ly�g��� l���BV�صi$az�a�̰Ư��Jg��;)bt�����<�R}c6�B���-;�2��O�Kc����PbO(o>8�<Ҳ��P�ӰH�2 ����#쩷wӱ��(�Ѡ��
���Nì,7�����B�۞k+W��I�!�'�����1aj�M>�����L��&��?�h�'>�g�,���J�����`nf����`��F�w����'UM��i�ߔM��������Yz�OoA�����4��Ȱ�`�4`�'R��3V4��T�/�6�����?]��=4t<����8o���~������!%�ڦ��CD�[��_<e���'�M��I̞���N��R�}�7�9��d���u�Yw謇�����A8	N�[����r���S$t�9�.3P�z�SZ�����1�(����Z��TAѥ[7��k`5pқ��@[��v�-K�G~-yyj�Exe��	eҧ��3e{~��:w!M�y=O���nl�-�8[���M��:�*���RY	0ܽ�V�DH����=<ќ�Z�F���ڶ�/E�Dc��
�]	�c���q�A2�j����6L����׼Ȑ�}�	��!T@��ʬh������VA�$��N�E�rf��gR�M�D�rI�ML�Y��dO�@HI���g���l�\���(�]��DkS��u*����)��%�%� P����V\�LF�HkZ�3EG�!ȸFĕ*j;���ō��HF�s�{����c��t^/�M+c��}�\�\"i��5yaX`7�';%[YfͲ�9%�Tj��x�f��V��u�K�퍅^��͆fA�F'��7���N�S�S�L'�[�׃�q�m�r\s/.�(�6��o�Hy_��hYIu1#f��#���(c-�2�kU��l^I}�ɒ& P ʴ�G6!�r%��׾��*7Bz�zC6\����r9TS�p}���c�yD���D>WXጟWd��d%T��ԓ�u�<����(�C��������]N���3� �B���@vƧ�X8�N�T�Ӆ_�"~X԰H���te��P)Ah`#v��C�[��%��j���|-��7���2��ށ,��{�W�,\�6���􎊸���sn:ݪ#Tn�A#I����n��BON���Dn y^�A����o)���7�*V%-�nx�q4�;�	 E��Q#��1���+d�|��O^� n��":1rQw��|Ґ?tH��l�Ni���W"����[ 7~��b�-�����"P><�{4E���_B���J�-�z�.#��U"f�z���q�����<bSN��Yꞿg`�����-�@��P��Rك�*]p��=e�ӒT�k	�A0�v���X�7�0ppZ�#B�>��qh!U���@z�ol�zb�}�G�s *}��qu^��b����P��]t>��M�
� {�M����[�a�5� ?���ZY�F�ډ��:�~D. :�q����v����i���f'�I�;��N����X��+��B@V�F�7�p�Ϭ��W'��~���ԟ�f�q��v3J�g�C�l�����k��X�#���9��n�\�`���
�~k�b�QuO�rq6O+zV녕��_�=@j���JS9��{�Ǉ�.�A�ب;�T)�\��H\��| EJ�ڷ�v���q��A�G���e���^�-a��WIϘ�`X3��
-Y�kK��13�QM4�Zk�)�W�S���o�h5:)�Kڦ[��C��?֑� �-���>�-!i��������C�(��W
Lp�~�/��S�0Yٝf^�(���A���[\���j��cj>Y�s�6U�A�h �谎T��p�x�@���NARu�������}��m}`�kj(ڀ�]R����`U<��	u�U��4��B� ��/�x����J.������V����o:��q�C��
��������卵a�%�/��YP/�V�D0��X{%��J�|��4�6�MH���l���++=<%�C癸��͖t�0V5��j��%y��QOb{���y����{�Nby?�[���ع��m淡?��
�B�Me�g�vvt ҉��ψf�6��4��`��@8�[���d	m���m����S�y�ذS�`�)E���s̾hkus�'4���I�U8V�l��^�����*�p���.p5�R;JT(����;	O]��>^<�8�)Ý�D�ɘ�c�� �=Z�S	��K��Mz�&�<i���斚{���b�F���<��ǀI�T���-n�8�e�� ���P�Z}Ɍ�D�<�f��/cqk�uy7Չ�'vOf��mK%����6�Ph���<t�P��û����>�r�J���w��yz�/�kD �e�21,���m�y7�b��E�b|���E��uTp���MX�1�S~/׺y��Y��|���*;m�b�X���	��[�B�x׎��Crfuٶ�^}Yr@�X��c�Q�T�l��\��5�
Κ\�ی��@OE�H��w,d!���PF�z����vj��N���7�g��"_�lH�� _y�V�yW��%�R�>�a��!�(Ar���0������!�
U2�O*���٫@���*dK�6�}���U�o��w|=!$��,���8�J�?s��Q$0�c��I_�Gw�d����8��:8�f�.��:�d ���W��!�A����I�g�dx#='�Op-	�çoE���!9���l��$Bs;rsg:�c�l�M�&�zy�.�t�U�|���	B k�j�u���v���;C9H�eR��<�<��B)ӱ��cJ�$s>�=���X�����\+���k����HCG�y������vw7�x v��T�/�'�&3��Yu�j���D����ɭ}�/�����Oͻ,�Q�d��Q�'!1�^��鄰|@c����k�G����G��(��ačA��#���?��t����Z>�1EBh���OXX`�=[�4rIk���ZJ6��S�2�[M���At��/q�@t���������*�������6`�Z����WWm����%Z��𭒼 Vn8 ]z�ρ�a�����;���ʩ�N	�&5��GDh0���ck�<�?���V�m��)��lI�PE�p�����e��؈h�Cf^ɞ�^��)�V� ����
�����ڕ	|*2'�6�����Q|}X7S9�z8�jqK!�����?)��e4C��ϊ������g�$��Q u�s��x+�����(��!�V�9d�L�ǈ*:qA�q�%�hc=�+�#���4��4��Kmv�0�ȷ_���s����qgV����A�,�su�h���6���=�����ȋ��3�ٿw��o$�J��r�WZ~wr���f���M�^�
�����]v�rߗ>�p�� -���1ΦGboq`�}M����Q����ŽPQ�YI� O��yO
���Ʌ�ٮ �	S$g`4"'Lg4���Γ�#{JC;.�~�>�/շT�
	
��s���ϓWπ�Y�<:���=?즋�D*��<��|�OX03�W��vO�P��l��L�;���f��H��ʼQ~v1���t���ݧa؞�:D4t�l���NQ��N�=�RNY&�����^c�G����[`�>���y�����6�3C�
8�*�YD�����)!�Q=�(�}c� }3�xb	���|�)�s8lz{J���l����)#��ȁ'՝6-X�|��)6�e��SWدG�*g��ˈ��E͂Ƨ�\��G\8�BRuUq��`� ����o�YĮ�Ծ�H����sO��*�C�����_+�9Qâ�9�z��@g�ڧă)���g;��c�.���h%���"�z�h���"�cq[�g[II�`|yd�Q�x��i�v�5�rQ48�(�S{8�D�X�A����F��n,]lc��c3qovbz��J��N�D�����L,F���KDN7����j�!VsGd�v��@ȤD��	���ܭ�1S��P��d�a=��C�B֤P��a/�.Tƍ޼��#!�^#z���3V�7rIt��2�pJ���rp��ǃVA}=��eԕ����ՍV;u�p�LҏS�6[[������Eb�X��+��L��JѲ��_��y8S�-μg�g+�/;^��4?Զo���hg9.`���"��u���5�G��gj]��N�
l��:�~ٴ���$	"TN�_���E8���%7�k1c�xTph�ִ��v��N��L��`a6��}֤{�������ԉ�����^�zn�ƛ���hdx������p��9�-�	Z��Ůɠ��Bm���m��G1�tצ����;��x�X���N��N}�o#Ep·�F��s~��
h��CFs4+}S����*Y�S��{_�^�I�����@wa+޸o�Ҿ�����eN������>��bUؘp9)�Ka���p��j �2,5֑�}z&ЭԐr�)8׿�gM&���HƂN�� �KX��R�||��~fy}{��>�K��vǎ�4���ҵ7"3v5�`��i�1�E9U�**I�y��w�Zhq�Q���$��pYk��7�̋������p?�D���g�u�l���'Eޠ�������0#,oj�>�p�M�Q���T j�ZF�����"��"�j��F����N�!�<Ͷ�a3�øh�BW�b{ƥ UA��!޸��m J�'5�d��؟ȂFz��w�e��Z�)�h��H�L$eef{W�Q^��e�EK�tA������
�x�sf�&A1�p��fQ����pT\�@��n)�?%(����n�R�r"�S&�y�+���.6~��CB��oY�-�n��,��U�տK����y@~���(�RP��b�����T/�"��i���#PEҙ�jj�^��F^$4a��=�l|�vZ�˙k���C���c(��1Ӽ=Q�UɃ�'��.*ޥ�S9?��k��]�H��!Z�#�1�F��֘e�u�W6˖�B��mf���OO���*7{����5%����g���4X��Xd���� 0��F8�5���4�&��[f�9Z"��G��y���H&ٺ^��䷠G������r�!^�F+�<���h	LS�\H.SJ�L9��ѐ9'[��p�������t#Õ��7��Y��1�AT�|�}�����a�7.6����zE�ml�_���j�Uزz�>���n)���*�ө	ϝ궷�_ާ��f���V�8����+�@Ȁ�0W��(�+��}~��`�F)��9Y��װ�l��Ӛ\Ðyi}S�$ھ\�ٕx�(}z�)B�~ɐ��)["UK�-�@/xL��}�֌�!Ճ`Ȩ	�>��g6�L}��۽��;��>@�&B,�/0��cr���_]�ǭʌ���a4N�Yx��h�'K���]i/I��@�7�V�a!A���)��l�<И�Jt7�~v�[A��ާ���V�5)p�|�8���Ö��0��r+�A���M�R0V]d��3#+�n4�.�}�s�y:����/���n"k��ţ@�l�y���?{`mh3̐F�J�3��3�+p�ώ��n��b��)~0��f��ճD���	�&��Y<[y z ]�dkc���K�_"���K
�jRKՙY�� ��,�Y��FY��T9��]�^�L�M�@Ȫ}7�k!��!�3�|S+����׌�3�n�a�X��_@d᪗L6Ym�^(���T�	P�'y�4LhX��A;br��S�]��sI���u����f弲bJ(X�h�K�G�v"̻�ߋe��V���4h�ƫ����K@Wq7��^�{��,�~񲘚uE�o��%d>,Nx;b�e����Z���Y]� 2lh���ر�X�Rm[�Fi��Rm�nV
3�������m;2%
���iZ0�8F
'Pei�n�N ���8E�0"����$�o�0B���og󛮯U[Ͳ�s���D)h5�v�8J��x���������lg3��\���F��M�C���W֋�� ?�sP��V�B{}�r�bw�d�ԒK�f@�.�LnC�f�1{Zqhͼ��o��C��_�M�w�MN�Ui��1��0Ñ{�j1ٞ�u�e�)�p�͊�.���ݶW�NW"/q&?U�H���
�����u�F����Kz�Z���%�*]N:�Y`��@����eQ�_�U��'��o��F�2�w���8��1�J�zz�y�����U���n�_�.�5L�I�-hP�C�������Z��vG�#��M^���&w|�|Һ��S���)�M*MF�}'|�\����q�����J)R��J�tk~(���3��� 	rv�9M�˂�a� i�&{����&5B慱�IPt|�*�b S� ���YV�Sh�f�!%S5�o�r������w�N��\�{SH�e���� 4��sÃ`�w��h9!�+�> ���������|*����s�<�K�ܒ�Mi!�<k�3��?D"����4�b��8W��Q�O[�9>�h���v��@g;L+ٛ�����g��U���Rֳyc��9JH ��b���q��`	���=)s�b�|��9�K��4��	�� ���?�nOC#=��� �gh{-^]���Qs,u��c�V4�
t�Ȩ�-��sӂ�/�x ���+���K�9�ϧ`�
hRȪ�Z��=9ɻ�v8�����%��{��Iњ�KUG�1�|?��k�b�N!����b�r���o�ͅ��e���0�Hki	I��G�iO_#�a͓�����K�>�p�.Q�_��;ƹL^˪l@��]5�@��x��?��W�Lg?Ʈ�9����.2m�9i�v�����=�<W��p\��ެX�f��W�\m� ��	���/��x�����u�LZB��닉�	�_Sv�8�m9Z���$z<�����x���\�/�e���n�e��6�Rr���d 6��B���"d@�t��Hh���<�6g�ʵ;��%�FQ0�Yts0�R�������F�򜍓�d���fyޯ���,��/.ŕ�u�s��^j�X�,�7ZI�~�8�)}�H{3�f��0�`�U�h��\M,��Q����i�f��{���>���*6;-U8F��j Yp�i��ա�x�@��RJ��"i}߁r	�r#Lv-��!%�&V��h����$��a�I{��V�e�� �9|��Y�t9G��d�g�V���p�Q������kFy��}�����WiXk݁�~#!��n\�3�*�M���9�
�Mӧ}ѳ�qt��v�ļ`��֫�	�a^��$-�A����6^I�`A��b$�K�T�
�q��Hs���3���� rZ��1��H�,`����~��gkZ'W""��ʃm4��29G���Y�L:�̩�7l�8*�YZD�?9�e<{�ފW������]j���n}�;�%��c�Zέ ��"iO��a|M��g+D�F{�`�`	���j�3��nu���l�,�0�q��H7�~�_�
΃��0�����W�<��\D�[�VU��C�%��1���.ȕi2��-8�ӧcl#���#~�
�U?;���ڻEW�w`�/���:ڷ~�9eDK��d���s|�,�q�{�	dQQ �W:/���	�jw�0�Kۭ����'z��^Ŷ�$��|Q�-�E|��Ԕ7��7<��&����[�Ӧ�R�5�:�4:�߰�Wb"e��� ˳�Baᨿ����5�@㒫}K4T$� ՚d�J��J�mE�W�o{�A?�A�=8Hq�w�C
�B�m���AV��=�
����b6ukklx�� [�����7��Cqv�����<�lʶ8���PU=�[e��sG��7F��\1h#lq��bܻ��b6c�Τֳ�_�w�s��r�lZ�aR�K:�G�`E��g����A�x��&?57q���������I��� M>A&&Rb��T�I���_�j��C���_Gd��l(ڥ����_#2	��4&�i�WS���pGD.���m�i��HE@aOw��EWƸm�9��6I�׷��S�c��杩w:PBdOA���R	)5�w�ÕE�����#&�����$�-��uav���J~N��;��2��-��W#�S{Ѕѝ�oE�"b�����c��'��P<�$�_����ׁ����i}�ڿ��)P�q���57Ґ��\Uh4���ߑ�A��h�hp��ƺ+�X�}���Iesң��"f=uw�G�s@�;�ղ6����D���0uL�̄52[���'��*�O.�y��l������p��!n��]�+*w
�K� `��܏��V<���e?�0I�����f�:8��o������߇���}���ɼ�5H@�d��f��pwlL+ ���C�+d�0��og�O�l��:��PZ�ČY#� qF]����6��O\2�J��e~BJUI�<]v@`Q�� �|̜N4B�ӈj?�H�!�6��U�z�9��Z�����*��3o5�ȣs�6!\�䪌����{'ƭ��4��.փV�Wަ���]�ǭݠ�F�E*!���a1�U�qK��[�:nu��[*��č^�=�X��(��3E���S�Lڱ�$���D���.G߯���(ο��ΰ_7t��V��ҡm�"LF(t�Y#P�@�%YI��&1���s����)A��'�P 	j���s���
��D)S��[&.��<J�b���ɾ�Q62f�[d[��u�/���>���ɨt�jXŞn���͜DX��CP��,oP�#�L�v�D˼��( x �mPڹs�Ἢ��])�|�ym1�!i��yq�����\[uN��}�����a�n\��Ɂ�V���6��@��bJdg^�ӣ1vz� � �$��5fbg���5���T�2��d�%��'C��T��(�1
t_ j�bJ�J*�͏�f!J�p-j�e�E���
Q��I�1�©4��4��r�)ui���{XT�&<S%u	�}X��%�@��^���O�	ƈoVD&�Э�A�}��TPrH{Ѵ�\Xo:�q=�`��M����(�'�4��1�~U�%��Q}1%5�_�i;+
�7���_������(p�|�옖�Ӻ/�֝i�:��-U�(�T]��f��a巎R�������c��%�L�N�Ԟ��`��y���|�h�qD޶x�-��"b9Z%�p��k.Fwz�x��b�����߱=>l�_�	���xT}�\��DgB{L���'Z"���=��ڛ�WH�+E�9��*)��i(:�w����rb�������^�䫍ߘx�&��r���������-�^�o�N�@h�$ʳ\����>�V�ܔ���|�T�=R��?�뀵�)M
���f�d��d-8�����&�1�=~I�����#9��u�7nPC�s\����zO�n��eh�Llc��F���_�����(�j9�� �h@R]��p7��^1 "���.���'�Y@J>F/<��M��ƚ��8Y�^�N �۴��Z�����G��w���~��m�F�r�:m�e��h����]-,���z_�/#��).�%�G�i�1�
��Dg �t�uG�^J�oHm<��q���؞�Ok̈́�$L�`�b�l�ϛ�n�҉�su�xخ�T���{p�"N}X�H��W�����mh�?�2#����u�������5I]�����J��������qSU��,�sv�=�^%fW~us���&�E��&��PG�Mo�K,�1k���m3�R�~�P 6��k�k(+�V�A�Rj\�Ml���[ ��})>���M��dp~A�ӳ�O\��!��b��2�ybi�x��F���v�mMEM>���Q�.��WӰ�00Xp(�u�e1�g�`Ǥi����&�������=�1CZ��}lA6��_��R���͐��+���Tw�<'͵�c��o�M'��Z]x�V�r�.ο����% Sz�C�1����4����[�5�Zԩ��� 2��IY/�\�3�q�@�l �Ki9;ψ,ܟ�o���"vȂ ��.'�u3mU���>�lOV�XD3�)�GT_^���e�R�0/wfoG??;BևS��Keb��ӄ�ܾ����o�?1�w�FBa��F;�C�O�TO=�7�^
�A�CM�`�tu�SF�0�		��g_R�w#XT���X��hG�q����`s�C��9D�/�H��F�\vR��%"=�2���T�	����즿�x�DQ�F&
��R��
���	��؂��:d0�f����ֻ|J�pEZN �����n��L�jd���8��3�.g�$�hO��(ŰW妚�1`� c�q�W�\!����w�xd��2V�Č_���4�����L���]1��~,����=+P*��e/}6�:���j�1DmԮ�	�p}ov�~��^F�n�t��F�ؤ��z�����5�[fo��g�ZY��Q���%팇
�쬁4�|`��]�>�t� 7��<oT	Y�Gf��iz��{��U��>��L;�17p;�H���0����eG��t0�{p��ZɺE�2:Ic�A'�+T �N&�4w��@c��SP����w��Ԑ��(�iԧ�H���4j'������o>O���d�Q�={؃s���������ϴ��k�:^7�d3��"��$h�o52Ͱ���̨u�z���_�z�y������<�rr��*z�����`��RR6�b��?�ߚ���s�K�'�j�/��g���	a���,��w��/%w���]�~�*�����!��%�^�q�F4��0t���{�"��� �[��t���y!�	e4<�k}%˶O\��!={�0+.��@U�2-ٜ%�*n+ު�Т���G�4�����v:q�,O rb����H�l"��,��V�9�Le�ŵ1�TM}�O�
���}�_L]��K�tI)�J �8�H4�O�0��ʉF"L����o�5S��5ON9��gQ@�5-�5)��@pA��y�/���r.�d�6$����q���ؒ{�)=C���� �jP�=yf� w�$ ���J�=����b���	�Q=)O
�͕�k)��d�?=��ʬ�?�:L�Z	�4�����,�E�hу�P��!&�9�A���*k�3���k�X��̓�&�Ԓ�ώ^2vu�fZƦvWoݔ4�LV[�4 �o�~%@�M&%�x�b�j!%vzJ��(aD2�-�kn����9+P+��3$qsL
{J)�#;�]3��R���3]�Y�{>���l���p�}��f��\����8�(d)���;�T��3Ȍ.��w~A�����~O�5_]�P�L�d|�Q5'A���@�j��Y�P�T�K���=�Sc�4W*D��&|>$a�H=(��wz��)��'S����!�Q��w�	ވ��J`J��kT�<R��S�b���Z��g-�m��5~�4��yZk�k�n
�s���;�#�=ƒ��� S�a���gR�0�d�����vˎ�R�/�q�x�`��B��D,��0ܫx^�ڽ#,�w�wq�(9u��r)�\��PA����BG�G��YuV�e�"r���=��[�LS�����^���R�>4�x5����f�0���t�q�*O��U9Zl���P�G�, ���ޚW�X��"��J��ź|�t�:��<Hϕ}��������K��V���Q���6����.0�Kj?�=����X[�՝��Y�ZI��4��w���cb}�a�v��=��j�Ֆ���7����Ȫ��6'!`�2�G�'s�vU�f^��)Um�����2�kC�m�y��G8�+VODw^� +k��.��;Ә\�8�	���_���p�6o�!ზ[u��(��{B����m<3��D�*���u��s�A��`�"%��h�����8C�.bh�og�AsmQL�D����zHs&��9ɧݬ��M#�w�[V+ϑ�\8`_�E�����"zh���6���Ѯ�wB�5�q=a�+Ղ��G50E?�i>N`���w/n+��b�#	6Y��*���Pб�4S�g�3x�*Rм9Cآ����a/�n���F��K�N�V9
�ˉ�H��\b�(j��H4��Q�Be	T�������{[H�~3���M�UC�Iv���
�㝷����Hߓ�c����� v���
�2;���Q�N �kq�!N ��G��ᒏ�ؼ���bP�U�=�gI��eul�_���N��U)z��q�;�F0}���R�!�l�$�j�3�t�)!�� ʡp��c�o�� �5⢟�U2����XEJ�}|��VN�g�9�s��=5�kLXۼ�'�I/��TIM���'9��Jg����V�	N/��4�pKX��[橖��S+b��Ǚ􈪋��N(��vr l�: $��T1G��(K9�� 
�\6~���2B&��d/�z�σ%5��[c��`wUT�%$)�}l�^�8k�>�g�2���D�*H!i_\n�&�Y[�r�Lx�M���݂�VB����ZFs]	F�>θ}XV}���)��(I��m��o��>�/~�u �y��]w����}ʉ#�����p's�Iҁ�ؼ��3>��ߺr�n�&�ņ��������5E�	���-=�>?�7�	R\R;N�7\/��ꝉ"4���H��:esA�w�k�|���!S��1R.���y��������MM׸	d0�XB��X�/�ru��۳B��S�ru��Z $>�f�.���sS�s��S�7�Ah�i_p;��3��Q��q@*�p�as{L���h9E���c��(g�$ڕ�N�ѳ���s|�;��C�{������� )���_)l^+`E!ʇ_������c<�E�͘˴KY��47��V��0_$�
ܦ|BF�{s��ǧg��(��L'�w�.�0/g��*�\�>�����H��)Y8�Ǣd�x�U?]�Dӭ�n;��f�ͩ[�G�����e��]�����2�fS�c�3V��|[#	����e���^�4��(;2��^�Î��%(X"5�@�>ͲE]͠v��\)q�W/Vjg#����6�lU��+;:(: �hҳV8����Lg��{��������1t�ca�j�fu��h�86]�HL���w��mJ��>�mS�m��$�ѫ�.�"1vԌC����9;Zc7���/yz�uX?[�C�"&��҈���e�a!�f��|�v�h���v�[[��t���Ua�o#���e���x�06G��<�R{���_1u}�Ǿ@�_!j�t3�p;���Ox��V`���;�D�㝝�3��:�o���X�bL��PL��P0�ao�u�n+#�臋օf�Ն\
��c�����-Q�w���c1;��
�(k3������C��? wŔ�'���<%�4t,�3�&���X7����7}�2�%��.c��.1��$st	hK��#OC\��7�b)D�gj�;V�@��:��Y���̺@���1�3������0�y�����}[qy�[S,�P� $),�y"�ݰ����Z�jW�0JS 4��gOm�����\迶 ԋ�ezЏUI�ԭ~¯��;�T<Qp�3��'<
����BK>�F��dEN�lvx����p�*4W+8�r�N�P��"���>IU���>P��7�V��[`~�&jh��@�&�`���$��uT�6�=N�uX�~�S`��Z�o4�\!�d>80�G�w�d9[ B!	GF��}�dy1n��jI��N}	x�'l��!���	{��V��,@��D��,aV��A޻�4j�V��3�J�%ٝ	�� �D���璠*T�*�5�u�w�z�wdܶ	�[�QC�RaP1�팃���M�ȳKEu�lP��q"� -#�{��}�G��6�Fz�ۺ]r�z�7,���[/r�X||' �_��R����_�6G��%KP>���3���*Y��w�3��[,�W?��5�mx�ߗ� �,�OS���x��������G�� ��"��8�Jd���5?�wQ���-Z�ڝ�2�D���<���)^;^���Xb��0L�C����](g`�2RY*����|G���s��m����>k��?#
Hj�q��`��q�Yt�L�Vt��gW���
�2D����Ԉ�c�A8�vFk��"aY�Q��+b������8��A����lԲYv	�E>�N�ǞKZ?�\���0U�&P��]�rX<����w�^5�2̗���lX��Q_�D�R�l����?�"̾A�:qZ�6�k@aGvI�~ݼ���h����Js5�C*�������x��o�� ��p3\������OנZztF��~���]Y�p^��kϹ>��nyL@�a��H_r�� ԗ\6�o��{�%�yI��kU���N�mH���m%���G��(�����R���'���@\n��$��� �Å9=_�)�A�=HdHs�5�叉��B�՜�.X��=��'�_N���*�~�{]�d�#�XuD�O�h��{�-�^���������ʂz��
�O���������U�����='N��"߳W�x��K���w�Q��I<�)�����5kL�XH߀���V��?$�x���8wa�	cS�����Q�9 �+�/���Or���mW�hq�u��-����
�_$_:&D�_�I��"O%��n���;�vUT�k#d��LN��3����r�쬒��y]�_�Ȟh�f�ɢ ��o�^ʝ��@G���/vD��NQ3YcFaa�n�����ȦIf*߬����&�(�<�\�df����
��z�Dɀ([]���v�9�#�`b�`ʹ
$3�GU�@q
:�`� 2��ŅɆ{�b '^�9��C�tLj���ݚ����@ 	[�➊ஜU?���8�!6:����a*/Ŭ"��} ��G̵x-y	H5������ `*�1������=�[��;����w���uj�6B��D�E�9���"g�����evP��4Q�m�-����!��� �>;�`;���}Ex�W�:�C�dл:$�&.�)�o=��V�5���d���p&?�Pt���O�Q�`�ԭ��#���|��X�).P�_���<&��p��[���3"W;�@��T�,�P^�ȨQ�~�\��[�q0�D��N�tr�t�Qrs!V�߷�檄h��ذzpt�ylz-2U�\Қ���|��`ꭅ�b�^h��A?�k���6��B���_*9M)��=R�oJ9,�m��ae����G�\ (��]���ܷ2��Ep�4p�cv�ߪ؅���^?i���"���CI�J��mw6g��:es
�AA`Tͅ
��xji!��o���ic�-�A@�a
�=�A��M7�����w�Qu���"�"��`��{b��5!AS(���ge{+_u��7%!���h��v�[���W�-�F(�$�����B��鈒g��Ҟ�(I����鱓�����?1�)����D�@��zܜbD���d�.�K�cu��v&a"�5��Ӓ��Mr����^�n35�s�/>,� r�1	!��{��!��ѰCfr~�d�(뵟�>�>&�߹$4���-�cZu�/��0U�$CKګ�������x�F�O���'�!g��K���z���_��9�}�[`��5��L����u߃�+=%��TǓ��2�e�M$���r��:�\B�{}A�q�ײ�n�����@�� �:S�94���x���B����)�[ҫLS'#qr��R�S;0�e|�1�«kg#ԑ~W�J �[������OG�A~͂��f��Jc��d�
���];)fd��Bx�sjM���r\;R.�w����4=|Mv���OaK��,@��3���& -���ޗ�kS��e�����D�n�1�v�P��t6Њi쉍�O��͋��Ts��.�.�]s��qN�G�����\��!��:�N��Y+
�y�Jj�UQ�����ȿϸfۘ���Y[�d	%a��&�b�+����T��L�l��eg�[1}<1Ǿʯ��m�Zr�����a��Tz̽��3
�`q*�m��L�D�!������ʘy�>HB�����FLv��lp@�<�)�u��o�&�R�
�j*��H�ݍQ *N/h��E,p�D����QI������ؤ���W�zu�۴*8�V��- �M�G��
Ob@��{���w�YT����aqqh�˒�S]Fӌ�zTMҐh<e��9��r]t�7��rg���^����w7���6��{����u��\�*J�Rl1d�+	�l��Ӎ��7#��O���=�sת���ޱ��C~�x�) �2����]�jx��JUĸ�y�n�V��@���>
sc�9�����6�h�ؐ��u�+���{7�B<�ߘi�-���C�U_/u@=���A��`�m�%��;��Ԕ�ٙ�Ra\��tX~�R�"K8�A�R�n{,���U&����k�=0_߿�2���g�f�|�Us����q���	:SR!���J���֑;�h$+5�p�H��ÚL���j&ށ�p����&������@Q���f20�zQ�-�s����$�ʻC�o�� �����|
�T���M��a,�$�`4ř�A�*�B�dB�"m_���i�*Y��pgn�=�׶8��L'�6e7.,�X��s�-4<FV㫊g���8�# �;�b���+�S�0&&��$�����s�$�V�rKg���J�8���]@��T~�a"Fl\"�/�yv2׵-���P ItS��Z�m��N9����iڠs:�6��j�Yk;?v�t�/�p��z#c�D��M����:�z��0�q��ٚ*����w�;)���	�wz}�һjQ�ڊ�"Ur77!Cl,w�W��`(?�A����B�u��v)F���w�惀O�UBջ�<�Ƅ	'y��)��<x��k�SNW�zvs�޲yD:�6��e�D϶<iڻZ;}�i��*��N�r��6��
׉��t�Ʈ�����0H�sso�5w�g�jŃ������E+I+~��H\2�zHt�!����d�h��C�N�T)b�u[����H��a�w��/��;�s^�y�i����������RC�>�v���7=BFAۥ��C�0+�����;x�+��Hog;5��>j>��7hͫ|�L@�o�"�"����Q LI�Mϊ$�7<r�'(H�5���t]a��H�B����_/�K3	-��+:W�����$�j�H��g%JjN8)�7��杅lQNF��y�'73����A/B�.ɻV������	vaۂdQ�#��==:|��e�xhzah��hl��h������%mP�����w���)���r^��Ɛ�-����K��M]$�䣶ԝ���4����y�ژ,�"v� ��� �F��ᐻ�2"�G�;�Pn嵚��q%*�Ė4�<��C��B>��'��p��I�i)�Wi�ۮqO�*
=�>�Xw;��cD��96��N���.r�QE�En�O�H�g���/�c�"�n���z���h�[n���<Zu8^+6��
sG&/"�
�GG�ƻ�-�Q|�Z9J�aQ����^RD80�L�M6{L��ٸ�C'Y-o�����`̫6�r���6d�t�d��Ԓ �Sv6K�1H-ҋ�D��#��^xC�^�r���q,�`�Eɮ�+�w����5���p:�{�R�2Ϳe����I3	u�sfRQ����nOQV�걱��F��\\�V�zK��b�홬iJlPWp!��8�.��u\-n���}pN�eZ-�B�tE&DsQ����sj�(��Ce%�7�9Ȫ�h��3ǽ�a:��BnZW����]�nq�"�O���t%SWX�[&��a,�Y��y1W>:�D�;�ˡ���;b�3*9�$}1հ�FgsvN�k����1H��ؒ�9+�z���/ĵ�h���W�ۛҢE��m��ڳ>�z��K�|^B��rqHq�A.a3�3��wEߺF���/�}/xi���W]}(x��
�z�b/�
w]1�l��M:��2FguF��o.�!�i��8���{}���]2�$S"G�o�̷#������fҌGz�cs�f��F����(� Ί싩����=\��9�.�V=A�&'��e#�kTZ�mK�V���:u>d�o9/4��hq-���~�g�ˀ�����7�`���� �UH�vS�A�"��ʌF�cU:BP"���\IL���?����_�t�eG+��Mf��'�Ɋ!�¸D(�g��%l��=۵�ߩ���qy�n�N���&8�����J��+�[U���7,�_�R��]:��GI�-��L[*(��,U%O������$s1��]xt��`J��%��y�|�C�2���3�'YU�hb�/*�M�i�uH�prbH��'p=�-�haW1���*v�k7�K(�9?�O�#x@H:rE���ƕ4r�D�*Oj��ь�QI��!K�y��qd�+�\����l_�'N����(�t2�����m4y�n�6�h]8F�=}N�P�������� '
'|C\�Yl�����"XE�cʻb#�`8?�^��(�I�{0�ͺ��>�J��G�]��tVi�9���J��D{/���f$�e�)X�'�{���>�G; �騌���t����7=,;u�A�K�7��(&��,�3?�u{�ܸ)�u3O�Oy 	�����7��R���O���=D�-��
}���E2�C���{e�CIKڵ��w�(�l�G��Y�Q�*#:Z�l��c����2JG��r���9Ӂ�!�8aV����[���oBŔ�ןs
�����~z<>	}�g�Q�,�>2��w.�C��]�������V��D�pZ˨�n��Ќ@僵����4�,��&p!|�)����#��}^�e�B�$ PBA��Dm9��|8�_����kx��c*�2��P{��@ſ�|>_�C r���Vp��6��p���m\M��x��c��fb+1䷒3˅���k�P��bE)�O2��������T����t�v����I?��$��i���"Л�Ɔ�[+,ௐ?a���?
4���F���%3μ+�h�?��h�0�s k�_�$)1ݝ�lA�8#A��
N����hצ�U0��~��&ŗ]�-R�Oc��O�/�� �J�&2IS>�k��C��9߂捠�qnd+�-�Y��L��� Ѧ7%0��~��=���|X�9���Ώ�&�7�%�A��BA���E�Lұy)5B�E(��,}�L)I5#����,����k�g!-�|�}`�D��ax��,}�U�J�;cr(�pWyK
��*A�|^��8B�m�7�O���	|��_(���%��FZq;��2_�xD{d��W���+%�0�5��~�ݣ]��F>h!�N_h���o�l�:���]|�\
cL5�b���4�m�\���n�����
(w�Ч�o�[�[+ m.H��"��JZ���3G9���� ԡ�v�J+�G%�r� '-�������z�ql/�ݾ��M���6��C��mJ�s�4��`�.q���� 7C�ER��e0k�L��Fo p�f�
*{�#�����u�,��m��y�t�3�ϝI�\��!���Ţ{��*u��Xd�=�N�Ǎ���ޞ�[�(��.�PA�j�v��4>��2�#���N@��&��b� 9���RF˪m�����M���B�+�`h���3� �Z�"���*�*�rFPS��S
�'T�F�]��-�U��C!�B��F'��x���.��	�@x>�X�PN��Sv�h�
]��|� ~	�cD�dq럆���y�U��M���`�������*m�a	����k�=�TF��G���u{;�,xR�c�5v.�t��-�%��_7ݨz9�P��2i*� �܊Nb��	�?���8�~��QV�;O�3�W���p0����B=��FU�AvS��׋ X.��|��Z��=ӽ��Z�`�'��k���X1f������;v;���c9zo��j�U}+u�2��z潟���(�ںPn�<��i�7Ȭ嶊��`�7��z��&��|���z|��:X���Z(É�r��H"_Ƀ�fͲ�� ��եsKVR���'0��E�C� ���~E|��b�t�k�^��7S1��D<��y�밹�IQ��
��~>T@`yf��mCS�C���,d"��> R�m{&1�������"j��ľ�`���U�{��G��:�^fLy�Kvh�3%ˬ\y2���@�+�ܜa��`��Dʟ��{[�F�0��?ӡ��8����J��P��jkH�W�F�z��
�3��3:��M�{yre�c��.8�r�M��)�RN�s�쥐�g�8��.E��9u�rql?��F��,���}�/�b�w/ZT=�m�#xR��N�_�(������`,.x��������[S�o���~�ؐ$`�W�W�1估�Jmׂ�a���ܹ�f�r���g\�����?��}s�x�-�	��CԦ�npf�~��Ȕ���>��a�� �|�2k����N�����s�h��͠�#�A=.�F~��@�}s%PA��\�;>sٿ DrTق�m=ۃ�i�Z��/�v�%۰1���h�/&�Y�	���Ds�C�\M�t핁Q��s���ry�q�2�6�R�ʥ=�>a�f�Dn4�a2Z�' ���o|��#X!�z��$��'���J�B�_�a\M򑰍�v�aKn6����6���}x�Eא��{�{���H�w@ɞk$���C�J��&dE_��Ƭ���u'H�D���Dp��>G�=I	� ���ܾx�ݢ�*0}�k�sw}7�W Xxn"�61<l��ܮay���D��������b
+o�d�3:�ݴ�%ֹ�*ML�}&�z��oY�gZ�n)W/�����PU������CEp��=�^�[ �7�?��/��j,L��j�:̓��@p�*�]����_���bu�\��[q]xC%^V��ܶk �[ƅ��� _�Tqe����)=͢��T��璼N�DY{o^fH"2ȇ�w2�g�ܚpi%�7e���'���łW� �Dl&2|��s�b�gWbTi��n˭=tX�_\)*������T�4Ho�VY�,�Vhc�����h��tH����Z�v1/^G&q/��	Ҹ�awl�9L�Z����A&��C�"����MUR����a�\h���6�� ��"��blgS: Ie����WjQ@ X���4���1Ğk�- �.~k*��U��+0��J�����Mv�o�W���՞S���EJ��4�F�9�3!�����J��t���AG%����	
��ݑ�z(��~������r��ύ`����y�y�>��I������I���ģ���@O����w�����	T�˴����H�Y�"��2
��R@_������Hk���!���R���B�M���#���)1�	�Nz�yu� O0yTQ��Y��LQ����r�$��ץ»���'�]hs��^�XI���q��Nɸ<��|���a����2c<�IpBѬ�s��z��5�"��%���٫w����U���uN����0�Y�}�����g�W�q�%�Cd��K��=��|���[������5o.��J(Z6�`��x�3��*�%�OIܲR4b�],f��=��BQ��JQυVFϜ��D��%�|��f�$�%����!�;����&�5Pof?���F{t]b��ʺ�T�R�D>���B'}��7�`���>�����[N�i���)�k�9'���RB%MX(��.y���*8¯B��j���.K9,	+_��+YҜP)��_>ps�v'����4����~��B�-�(5?���{.	���κT�c9I�g	�JooO���NQpb����e)�Q� �oY�/u���c�f��ڹ�%�4�k�R̲���Q 똊��9K6J0��7��A7����)+����<b��=�}���ȧ�bڐ����S�/�2��j�Q���4Duj,ʽ���I߹�ruS�ߠ�m �
�}J�F �����ۼ[�9������w�4�#���箇v'��b��8��|祗sJ)<lv���Ө��_�0B�(�z���	��QO�36���C,:o��3�x#�
��v8�|��v&�dŘ	̧�m���ħ��	0���L��	�f3�Ctu��G�E>�K��f6�o>I�	�`�5!,�Άt�DM)�����j�y3([�l�r7�e���|��;�2����+�\�ܞ��7@��4�4l���4��@g%i��5�Q��$�G��ޠ2�w�.N>��	�ˣ�'Զ�S5L)���!�y'��K����Ύ5���ZBӈ$xB��׳r�>���\�Eiܦ�:�ږ��^ۇ~���J�;�{;=)#0�xj�����6#]�E7^��L�}���@�a�Zf�櫹g��F;/g4��z�[z�T��2Z�H�A^��PV��J�v�y�e�`th�aJV���,��4G!��U"�C��溤�'	�� 4'sv���J㠡VR��_�B���O�)Y ���Sr��- �	��g���Ʋ�{ȭ�>�ǥ ���^�?�F^��x�&��e���y |`5�o��%���W��}���u��L%�\������G�9����|]�[�d�ѡ�Ƌ�`��Q�T��%���sQT�3�|u��B��3�ʭ��ђ�|w^B�^�_��1�o�`4���l�U�qQ��j��j�^�ϻc���χ���s��=ώ[=b}�	�5������~~��3#rtE��Z����Kv��#_�8#2m:�#�p�.M��J}��B�Y���̨!�ΏY Ā`&��AF�ζ@S�=�t��Uc��`v���CE���-�*��7Ps�KD�Wk���2��ͧ�`��b}����5�nf�5c�۔��~��h��vB%�u�Z��*�=�2�K=��Wa�����M������	���ͽ��6y��~6X���ٿ���tد���N@1�J�*���� d�E���Z�C����Ē�nD�`A�"�E��@!*���`TR�1�r~�+ ��f����_�v��PG7Ճ���I9��h�"�)�	��f�����������]�	�A-��4���F��.��'Z�Y&�L���Ёy�Ǐ�[��9�3�v��W�3�ˀ�Slk��	�)���4���v�!�$���t�C+ք1��L�ȯf1~���v��/l�'�`���G�E�X��QG��� ��ԑ�[뉃�`S@�n��v�k�p!u�I�K�%P1�5M��M/j�~{$��-Fr߸�il\���"�2{�\��lxQV6�+}��$j[*����Z�w[����I�V�O��5�޿L�^��*^�X���8�=�%Yd�u�mg?��Ǟv
5���L:؜�D;�d�kW���x&=�4��G`�}�� ��O����G��i�iI�B����T�5:�޾D�{��ؗb�������ꬨD,�F� ?�V������ۦ�J*Ԋ�G�N�5�]�yO3��4O�1f`���C6E���ى"fvs�^�m0M�"�"O�JiM4,�O��k��t� ��B�`��q����gH��ܧQ/�٨�Ȫ��N��YUe�!ʜ`[�S֝��V�,�B��(\H?
�K&3��͙T��)�_�)���k�-�kغA:a�+�nWr�u�)L�V���ZQ\���7���L�=pŰ�q5�^�3��a7˃X� ��1\�{O�ӈ3�)Ƒ��eW���Y~���0؊-�u�z!=��M�K�r�]d�k�tm������n��+Ra�9�Ǹ&��s5�_
Zt%���S?Y�y��rKq�2�����iR8Dk�b&����_�x��I���;�X�Z���5C�#!�Q����V���rN�ЂaC��?&�s�#$ƣb��a;5�<`9+OpE\i˳2W\8����ݺ�-z���K!�q���w<lC�RB�l�"y�2s��X���5�3�Xug�;��'	%��d�LX��)�����Bf
��AE�Bh��E!�����܃��Iڎ۾7��O��,��!.�㿏�㞽,G0現�Ef2����[�|�� ��/�CV�Q�l���N��I�S;@sa�l��=�S�XS��O��f���q m�W��:�ɖ��F���ZεpE3xQ1�5�6ΰ�R�W�"��BC�s5=ˁ8M"�Qrӻ �o͖Z�}����T"�.�xI��-`z� J�9���Q[�i�J��Ik6T�5�g��̒7����6	c���T�]���J%���e�:j>Wڏ/#S��FZ�ʤ'�巡��q0z�U�0c~v�K�iw�`�!����}�tq�]Էd�{��&�V�dHH,���Y/�)	%�w-L��E��#�d���A�,\�B �08�k#L���`��ت��w3�]�(�����;�J��9&uK9�
�\�0�v�hRAҳxkH����Z���8{��(��X�22����K�%@��B��A���Y�� ���ػs�h�m����O��C��U�&�#-C*�"�/�P��&���:�d v��a�*���:�(
�b_�.v���):<��u"Z�\���+)v��Xt=�
��[��T�e�O�P����Wn��u�ޑ��[�+l`l��V���v�i$�o�����ճ���>�wQft�7��a�mM�9+�s%���\�d�F�\uO45���>��@��6o4@/�jf��r4k��_��E��ʗ_�o����^2���w��k�<wג� g#+�3S`��<��g���x&��4Q���疜�v�����L?^ى�{`ؤ
��+����U�
.fC�7���{8�p���F>t�|T��=C.�� �+�]�yK�us|�(&TwN�kȩ�u?'�YR���b>
j��"W&���cv��_��a�
[�W���[H����b	���Q���@�sp�}�ś&f �Y�Z�X���X*�L�����͡3$�c�1�*�xp.�kۢkc�'�J
"�bu]00�B��Ē�� {�7|h��Y~��^oݙ�>]PT�=�J#��ǉx�?�K�W���+b�?�E��ɩ���+��έ�R�ј�:�5�YX��8�r3��i4��O{��"4�/������sΖ�/k�L|�P�>V��FA��ޔ�}��1�괮@d�2j�I	@W�_m�n,nb9��e2%���P^�����̺dd����C �y�u[Tz+%�v�_����7`��b�T�l�c�L������A�P_&�5���.��.-�<oO� z��=q3;av Ҁ6�G/M��}���8���ś���A�P~�)�z�����t���_w�z����c*j [��TN�Mn���F5�R@�Ndf�·Z�E��T}�}SEl��)^N���4�TL�9㕝��3�V���mY0/W�Ɋ/�}�q<kJIH�钿����X��`�|�mi�x�yQ%��6𝍣���_��;���eNֲ�>5xD&\��&:5����p�	_���/�N��U7�}z-ϳ����A��6<���'V�s2��3	.��3�8�=��	���$y�l"nl�9Lzo`�[���*���m�F
�좙hi����"�qi5����OQ/mcg�M���e��/O�}WY�v�>=�E��m���_K<��~��`�5����ן�J�^ʥ"�qQǳ�N:�;0|���D>R>!����Pr^�K_�N���1�Ӆ.����%��j��}�6�� �񞭟#�2�[~l�S����eviI�w���F]'Σ`���/b�%�;S��?Y���i�4�f̛�<��S�h�D����v���z�m�^6��FI0;	����0����Q�у(�T�}�'���O�E�zX��C'o��ڛ�H���
H�]q���:,g��Z��a0���|g��G�m͖���[Y� ���!���h��q̟ɞ�Bd���'yE�*�R�P��}O'�E�/�BZА_�~|���@9ϡ�1��z�1�~ӆ����߉�bA��brV#���Ww�	u�h�U#�!��x�w�* �:��ŗR�8B���Ͼ�W�8�s��T�!�f[�O����z������C��%�ωeQ>Y��4�'���\�MV1�Y즤*Ԛ�L��(�Z7�&S����G��P���ض)���dMFԊ?�KC}�3�v�h��U��t�*O���t��ݧX�7s�&t�Hp�P#�`�Z�w���dTf[�o��u�,X7������
d�H&i-i$d����\��.�U�D�t�	�w�$nn�W�x���-�M.�����n�vP��:���']��n_$+�� Dgҁ�W׊�O�h�.յ��Gco>"���+F�I�i7w=���)�&{J4n����yV���9M���g�e�*3��dϭ	}'5�[�'\^�ݬo\�C3O�rxe?X?�ڲ�o��j?Բ
��SW�F�X\��r�Q�xO���ت�*��~J��v�m��u�U�x%aT� /p�Ӽ�s.JTc�ĵ�� ǡ˵���B�����#1IGR�q-?o���S�7�A�<�����Y�pC��F9�8�ߢ�XI	$[���:<A�~�.�eE���.��Yo҄������ҡ����S��N��p`�o���i�4otn�@�J��l��9_�ݱ��9yq�ކ-/k>s7i]� /ӷ4l�{f�%�\C*ͧM���W�D��r+�?�}]�-y�@[�]��|�g<U�=_�i�/����Uƹw��轋��
�a16T�=ubĭ�a��@'M���f~�K`�o@�d��q�/�8� Nh��[$D� $����j���Q3hڛ���ZUc2іË"1������q`�Yy��h��^��j@n����6��Y�+n��Ņ~M���� �WV�Ԝ�/>�T��0�a|���g'=�ʉ��Xb�	��-�����]�b��wl!�N��q�V�6/�ۢ�G�A����j�R3���%Z� E:���¾���(ڷ���7�t�:�ٓ��bt̕�P�i�~5�䲁���Ml��4Yp�����=��$�^N"�u��#�۾�R���CtK@����f�x�ی� Zn��(�
�D�'�(���
��X3��/��8�O�|�� <&LYzn|U��k�]�"{ɫ�	���	JB}�-!��d��|#���H� �Y�����u��j�����X`eHsy�?�znZS\��t���g-Ǔ�<t*&�_�>�>�7�H ���(�EWU���G�#��A11�Eg�cX��ǫCYO���ҋ�Z�s����>lqP����C�pr�7$$�9W��_�#�F��H�7�役'����c��� �{8a����f�ztU�R#2$5'�4�%qyEb"��]�6FֻZ#.1�=)]�o� �~Њ:��\h?tY|�/@\�ܨ��+ܫ�0]��D�~�<-'��� N�/��r"� gC�҄����v��V:�m�{)u:�%� r0���G��O����E���_����M	�Ƃ������G��9
^�`�Eg�+�@~*o�T����'C�����sؓ�\��}T6�̛��r��r�@�wvB�crgʡ"��7�}�SU
&����f���*��x8�s�G����f BL&��'��U^\��cu�ba����o4 �ӭ�[���]������C�$��e�H�����?T����(�Sim�D�NP7�ô��-f`�0<�M9a���~:?�\y�j�ż��h/�:Q�$ �GF��!�f�c��7��� ���K5l7J	@���?�̛/T_-�M�Y���?�'���QT�쪰�S�*�i��$���~Ȏ�e[`�`�f� M7�7���z5̈́R�6(�/�;�gԷ��kGm���v�'l��M~jA�å�6��ˉjr����_t�^�7��q�{�w(��au!�[w��C?�g�I&�0��8��&��M��|�}���#:�L1�t�d�%��q�WS钻�Xq�F���1��h�U)d1�s��F����i���0��o�`D+I8�/Q|<��Y;�<b�0�8?v�m��<����B������"�lG��lB�[�TBȞG����ݸC� ���w<�9ߒ� �>����]�v�f�#J�L�_9~��8.����K.�%��@s�l%4�QI#iG|ieep�w���cB�w[�Z�������A��1��[����C��b�.�`A4%�Ɏq_d[����$���mS4)�w[�k�ZF^��IA��"E��:�y���S��߳����ͫ",�m�}D���a���/�gq=��4A�F�8e�iN�}6���Mx���2ǆ�O����]s���榫��c�@rV�iQׯBJ�n���]�>��2��������^��K�l^D3�]Ey��4M��9;�p�}3��m�����[�æb+w	S�#���y�kcQ �Z�3bVP_�>�7��� o�"�x��7�+T_���z0xs�mXɂ�m�
A%־�����+�W<�im�$0�Ń�4b~�ƊIP�Uq8R7.��M%�;�%b�OU�$��P��� `�uFFR1$�fm��/!XӨ&LD9��s�\aW(��k!n�̼`0��*#o@��b7o�^|o����f^H�N_+3��mO������?�ם���
np�^�^��wy��)8�0͇Ȉhf�ԉ��2��XJ�/�K�'���*F�6�l�gW{�ڱ�nq{�ӂO�ѥ����s_Ch@$��s
aZ�x�,"pf��iP�=�>3�x��Ҧ�Ц�o$vB@
T0	��

�׮�e��l.�ٲW/5Ufs�8B�L����&�G���qG��̷ r�K�G��q"X�H�u�w����<��Q��/̖��
SPq�����$��A�_3��*bL�ٮ*� !�TG�!��N'�Q%��fy�ŚR�S��t�8�n�K��Pa�N�U$�9�T��8�JP��J+�y�(e�Ap/���w�]'�����^}��4VY΁�X��C���s��ηg�V8�b�M�]��$N�b�����6�7�$'�+�[E�.](@A���K��%���������?�����7�]����~�&�U}ٿj��R�W{C�[S!��E�������{��������]�XY��,��n5�]���PL�V�E�$���'�@���2�Eۑh5��)Ġ�0	X��8U���t���M��2��O� �K�؁���֑uZ��,�u2G�����b��f�Ba-Q���0Q4�$F|��/Q l`�K,�!_A�đ��x�l_{P�x���A7���߷�&�.���)�:��bs
2���J4�+wq��b�ָ?�K�h��+�hn�E��Sg<�;GyEf�M���r޼o�}����3�g�����r,A�`,oO&���@��F�e�I���#���1RCO�|mbq�<�i$(�e��P�?1�F���E���
�p�Y(Q-��Q�̇L�5f��Y���� [
�������Y5�%'��{c���ET�,�R�=*�G5�=@��B	�'~��mHv59!�T�ఐur`���͸v꧄z�7�R�+&�T�MݎN1)?g`E�t����*�k��X_V�cvSXU~������2��W*�m�Έ�-�4�ٵJ����Y�1Y���̴	rC��{����v�j�T��ZE�iJ�X$g%���1�T��E�h�z���s8W�R1�>�{o��ٮ?e��츥���Mx�΀�,t�Cj�݈Z���DU��C��|�<0-�I^"��s���Cr�CG$U��c+�h��H�hT��Oa��q0���`�E1�}I=�!�\]n#&��zx�Kq�S'Ě���M�a}������>r��6������'\~�r@O�P��.)+�}�Kܙ>�
��rBZ+٪�=��r}.2�CB|Δ��`Ȃ���g���]���i[[�����fY�����~9�B�;~q��?Y;�%�����uc�Z�)���͘�(kMح��(���-����/��S���ߜ�
�q ���]�o9�U9ve?O���m7�i���
��'��:�{p�/|m�,/"H"���X��ī��K4��4D���G�w�����ֳ��-`�|����ei�@I�S�Lx�Ɖ�(�k�za�!�]�d��5��%�͔����%�3�����fc�*�O�<��c���!��`���U%!_�,C�o�@��ﷳ�jA<��n.YB�c�0C#��t}U�ǜr(���<��-�W$�QP��S�
!�Y�;gyn�.���f���u�W��c<J�h�e�>dU>&IT��t-�Yb��	���N��+����v���Q����4$���uTP�$y��?�Y�}��)2�����-�`	|������(U�U�]�zG��6�~�1vxlg����C�A5���*.@ۊ0�����ŋų�ˇ���P�o�I��( .�
��P�q�+��t�F'��j����ݞ|���B��r
f\���L?����ѿ�[M;\ni�z�R�'T�49of���؇` �I���!�.���U�#��y�ᯫ��tO�_�U�v\����0D�h��8(�o�)y��:[
��5��p���M��{��bJ!:ض��7l�A������`5�1�\%U H�k���Pj3&Z�8CD�J��T3�|?�ޑ6������8�R�8G쫠%�J��O����YO_�h��F��I����;�K���گ�X�����0*��ڄ2�~�	.��K��s��'f��Y�-��
;�̣W���
��X��$YZ�}�����C���r��g|�GZ>&ꘔ���^�Y�����Yf.�N�($HEƃ_{�;����T��%�����!�ްf�x��y�����k&���M5^Zqz��z��^�SX^3=E'P�=0f��ze)����A��v��|z!���'�]�gN��|�\)��g��Sn$��p���|W	e�Bx��9 �ވ��Om<V��1mڋYY�NK�|E�l�r�a�]Љ�e�(������9�I 4wGy�+�pC�óy���w������uм��rƱ�8���a��� 5�;(�]DvS�Z��6d�$#� K�� �1˗ͪ�;-��$�3g
�^�Z`�+`W!���7��)��\Z��C�Z����{�����fX`C�Z���U�iL�٣>��RKٖ*=�	��h�5���9�l�Ȳ��e���NI�%�r
"#u:�)%�3g����3���_���Rl�M����V'��x�Yu�(Jo�X���}��������Q(��m1/ζ�m�/�hT�����`i��65�e�"L.ƐZ_!�rE֝ayba�@W��)��R���ȟ���(c5���Ʌ/1�B�d�8�e���N��er��j0 1-t���}g�)� pX�|D��������ʛ�{_j�o��ƂR��K(;2rA�YF�1%��P��M���尗
d�ƙ����zxxjpF;�VB��I���;V���%��Q�\'*�������O����c�޷��($�Io���2jYa[ :�
��?��t�(�Ǩ�0����Z�gR7@��떗���'�,d�bxK��^#V�a~��;�@�}�3�L��3�i��C�DOc���,�0oԦN8\������-9��ZF�a��[\�#cӗ���qP������1cH�@��<��4�w����Z��a�hdt�p�1b��+dQ_&{���c�E�R�a�܋�N�?զ�Ӌd��+�8~,�s�KC-<�8G?H��~�@�EH�	�Xow�-v�����1�BR�w�!�T���G���*���@/k�K�����Q�M�> �*	�@L{*�(���|1�8M�gX@�D0�Q	�sQ4�q��ųb�B�RqH�>�Q��q���� �J���c�-����#:۟��tF�\U ��J��m����T��`�3�Tk}��� Y��qi���Jsz�Mr�Q��RW#��hs��ޖ<W�Y�� �]�ǳ�Fgt���
#��D}�M<�I�g�y*Z� ���-�a5�z7	t:�t��_����Û����{���wc	�m����ܷM	ǘ7[��oL%�ȷ.����A�, �u�������������H���tS��H��c�FG4M���8�z���򘍸I���H�$.v����=h��[40�##2�T~M���[k�kqL+�!�H��ċ��oE���B��:L���1�(��J\~�Z��K�P���-� �$~�nΖ��y��O�{�bڰ�s�b(�1���W��v8F��fT\��Doe�%�1D�qv��D�K�
P[�O�^g5��.�p�
��H��:{zI^�����p�l�5��z�7�.!k��K&�$�.�?.}n�r����͓ "�*�:E%�:��Fsӧҫ�����lP���m�zҒ�7fvJz��$]�
J(Ǒ��%,k�ݸ�&�R�ci5��
�[2��@m:��v���ŒTj�T�Q�fʹ�-ǔɉ/[��$
.[�7}�Z��s~k�A�c�Ճ���5�k]�5H�(���n��h�N�,�R/mCVZ����N�u@J�|x����£�*22�?k�Τ̉@�$�cޑ�hE��^�؏c��y�6��!�=0U��Cv	��/	�Vt*�S���z�ٚD3B.�JZ$&Gi�Y>Ԡ���a�K�H��eZxx�jG_�� ,x��dT�@B�o�'�T{˜P��][�{��×�����ū�o3[�P����#�0C�m�i�͋˖�r��}���Y���tq����ڗ; �v��<�bV
�\	���u#�ŏHÑH<���[�O8�W�n����O�yAc��(�C�Xg4I�y'�&B���D���i�*���)�k�ν��$2�M�P�D���O��+��yٜ�q]g��]�d�H����T��"���)g,b�z�'�_��U���|A�C��:zE#��Su$���_S1��;c���e\D�As��k 7�`b��K�I��,��(���$�[��|,��}t��Ó���Hz���[���T������Eו�&�;�/H�Ӎ?�����> �����>o!�N4Jn���3n�0�K$u�3�i�N��49z�/=t����i�˓>e��V�^�������<��'A��B�w�<6
�\���/)B�Q�= ���G�DԘ��[ֶ���&mܶ�>(H�c��Jȥ�^rfػC}fZ�1�ϒL#�7��������B���N�S�F���$�g�?p6k�W`T�a�!U��d�ON��q�cl����:"�
w���pJ\��@��`Qba�u]�#�ŧ٘��C���}��YZ� +z�C�PV`"3.07m\��t'e�K�6���Ɔ���D�X)�
̏q+O�U�U���ֵ��)ٍ�<�Xc��Ns[��^��т����HH)���)�,�2�R�+\�lt����g�dMԾ)Ό�������GF��0m�A��_q�!m4��wd@|[����s�0?����7)\�[�*$r�ܣ����e��C����^�ᒄhZ׽�9dm:_�{'m3<�~}���0�/]�y~3o��MI�
@�O��d�P&�h��wQB'��PJĜxdc���4 ��Ӻ���R7Hj�$��y���*��Y��Z��G��L#�?�BL��w���:(��#J�<�Z8����	�lKb�v4��K4�|��	��.|,��i*��P|����,sR&v��*E��Xג�E��GI^M�B�jж�G>��-҇G7�@F��������v�D����`�g3IsBk��KzjbM�/��\{�H�՗�.��?���T����V	�p�nE�G��� �׃?��t�*�Cs�$D�&�p�/��f�5J����_N1��i$^ٚ��g'n!~ȥ� �������>�tM�'�F:�ס>�ro9y���/@j��|\�/w�g&��-o�]k"�Ը��i�j�����z��ٲ�)HGv�1ӳ}<�2��ݶ�ȣ)����U�+{o�e'k�Z[�I�R�ޗЉ�h��*U����<=s�V��H�v�3�EKc��� ����[�*��:��|���I#Ӡ��W�߻��|,6o𩀘-Sv�"����ū������'�/�`�6��HfQ8t핒>�����q��f0}q��_���um�@�x�G-:V�6c
�4}q�%�x��p/�[��5<ٮ����%���'U��9�n���A���C��j�R��c��^3h��/ze�Q��Pzk���U�j��n��[5c�<Xɜ���4�#صШ"���ZI3P�Q`��W[5�wɔDY���@i�?8���=�B�8O1��
�z5� ��jt����P���<�+Mz�bE�DEĊ�s�S�>|�k�"(]	�q�Ԭ��U��@8O�.�mwr�-����1ZM��yk�����!����[7?<�&H�����>N�Z�(�;E�I���
�w��>���������F���Ko��(N�𮵁r�ĳ��6o�bs9$	s}���}���[�0�Q�Դ��lP�|z�����HM�����
<CFVMM*'@�O��c����f�P���<�Hn�����Ѝ�2F�Q�a�M����'I�}�k��*LS���k�/<�A̫�55��~�Lv��&���6C%&�ϖ2gȯ�$¢x�O]���&��i �E����Ս����!��:r�`���.:��a-���|Ȱ	gA�y켈!�>CR�*����j�Y�˨)�:���Ӳ./�sN3x�7�5 	oR���7��0|&�3�(��ɷ�*�����ʱlB��ਿ.� 9P��Y�i+By�ʱ�B%���H����UC�F�|� �(�:a�Yo���K�wi��=���T��,R��0j��W0�{{�C��^�n�\�d���E�PLұ+�i��*$#{�#j�p?�����u�_���c=�Ʉ
��R�C0O����-�-W���6Z�V���C�?�^���)�~�E��Qձ����G��/q������雁Ho9,-�ͯ��8��9D�>C�D,eyr(�mjZtX`���o�pت��#d��<����TW�*
gl����2گ;��6�]o6�
tQ0z�єR~z]��+�m#������8��ě�����@�MJj~ߎ�Iv��؈��BO�E�랹g�c7�G?{�D+SK�V�������|؊�#4����L�d��T��i� ��􈖧:�>��s/�f=ZԖ��͉��#o��x�C�<�?ܥ�쁨�`l
�jQ�m��{ү
Y)���-E��)V�I쑋��)v&��S��n�5= Ɩ��;t�-́��t�1���޼��e���![/��H��K� �߸�A�wJ$c���~�bF�{���~w�|N:����6�޳�Z�!�A̘�n��L��O�l�yq�i��Z~��@��3u	x�d�(n_m_��V��!8���1(rձS`B�E�#��i��g�����Os$�'�'�D8�?���8�&&UR�Ц� 
+�b�7�L4��e�H\̢M��!�s�Ex�=�"n�jHA�J�u�x�R��@n�No��^h�l�F@\������T�����L�CtP�S}�e�$��TeѺ�E�>�	Z�#0^]8��U��	I�$����e���X"�K�;y��� ʂ��2����I��bEv�>��/���R��hm�ΘT�A���:�(}�:lgE�R+��Pdu�CzX��6��pn9�~�ĮL�oj��^�����t��w~�c�j�ZYFi�+�U�������[X#�j*��!�i|�<��]���ϰq�JBٖ���L��kh�5�i˺�S&�
�a߉$AV�L�M�&�n��?�4&��{�A��J�H�{ϖ0
�xf�b��r���W���)��jO�B������`J"����*�P�lN��i~��r&�K�+�E3+_$Sڙ��&K��ܤ���U�7���<�2�Az9��I?]�f,9i�q��n�ڮ�""�2���68�������2>։����Kn{�5�]H8y�ξ�`������M@F��]D�jVH�A;��M�X+�r���H�q
��� �C}g6�kA���}�b�D�5a�Qk�1�(8�+���*N>�z�ah�g�"�|-���m�#�����>�/��IkҨ���.�]���r��7l�%;��!�}�����Ӷ����$��&ʛ-��Z�Q��WO�eD_���v�������Z�^�V7Թ�)8(�V�x'�{�ǌ�l$����v�d�~�+�s�d�C�&2�,LbȢ\3G��H����%I���PɁ���'�|�ꢰ4�m�xl!���ͬ������B,�_'�L��:�Ւ ���Hc����O�#1�`ٳ�E�2`g���o�ϔ�)m*��AB�
_�Fc��{
Rh���R�$ڴ����� N�;�q��n�F��b˄y/������/�a�y}(�`���M�\�T�x�IR��l��S*��g#dF�����{��?P��&y��C���� <T�vD:����W�;�85�4m�����3����[�n+�! ��#��SE�`�5�S>��V@�ݸ��WX1��+�0��#��և!����R\��A��i�{	���
V���vBKx��"؅��b�<]W�j��'�+�Ek�Mꑃ¢kqͲ��M8q�Fd�M,�?�STO�����Cl�`
H]��L\?U�;fy����?��%]����k2�{u�}�F�_��nմS�Hhh����$������W��c5�l���A����Q��m�!���?f=�����/W�WN��ݵ Ǹǅ���{��Sm�7���7z�ژ,��L�	�i�T��t��������9m+��^��^c��z�]Y�፮��܀������c�)3��z�<}ĔR��񫰏���FV�'!���D��>y0�޻�O��-�k��1���ٝ��4��9����)�y��U&���r�l��i�A��0-���]uE�����/"��8�l�\�o��;oW6H�u?-�m"&8|��d�����@[��vWq�z�c���8��7ǚK�|���x�(/����1"nEG�}|�/����-Jߞ��S��Ux��>R<��������c���"�:7|���C0���Փ�2�M(�:��Y6���H��P1�1��2=��r��m�	���R��uJ�>k�Ǜװ������pb�����@q�?�e��D��)��*t�Б`D	���� �Bj�q�j�C��P�ry��d���=f	����+�	^���sRݢ��D;>uіT�ϰ���y3`����}���߮kBN�O��{!��6����|,���hl/T��f_��"G���w�<�J8u|~tW��	���U=@�7\�꯸X%�Z���\瓸�:_�!�{�b���';,ݓ�&>$���1�{>��E� 39�g��e.��
������_#Zv�v��uP��,�=Q�7m�ٗ�t�_:���)�Z��'篡*v��+�߀q�e��-3f��i��y�(�I�e�o��O�۝Y�J�҅.�*;<(��^[\
I�'�V;��ʌY�Ϟ��?��|'-�;�K�?�@m9�
�}�����<�]��moD�ҳ�u�{R�zKӨ�AWu�
��&t)1��޻����V���}�]����x�$�9gE)o[�R(��S<�1����R)z[Ro��$�f�Dj�v�V,�*f��5��㑛��9��/�w#���B1~\������L^�PZ:�y+�Z��v�}�|j/�������\�z��%�m=��fN0��2I�����gc��L��>��<��B�����5V۽pN���5��
�����㿳B|{�S�j�=5���>�Z�	� �S��Ҕ�{r 4�xeʫ7�~��q�x#Z٠~v3�z��dJ+4w����<�7���ޅ4��@�{�%��ȉ��se{a��,\��.�A0F�I"	®�k���!5��z~�N���w���ֿ�KO���f)T������(b�q�<��O�f�ټ�A+4�`5�1�A�F�!��LX����5cb)�M�X;��#[6�	�X�P���8-�2��N������e�go��?5��E����'z��uu~��5tP�l������+Z�!i����j��dƹ=��x�!M�`��<���Kn�M�#���V��w���~��FY�i�L:��m[�S�Z�I��iw4�����\�+[��}\AJɝM3�+�|5�>*݃L�T=X�&������.���"��m%ؗ_��%�O쌉�͈���/m�����[����=�f�	4��+AW�/����&>�����Mt�ipo_M�W�@�46��t�"N��:f����DѨu�@���}����Jhr��5�����]3K����v�$9�e4QnԬ߰w����$z�vR�or5Dd#a<�nƅg�ʩ����_fL �ߐ�nC�Ik���+���]��d�� �}J�x�J��a�(L�]!A��\!ƽA��$�EY�J�Y]a�#�p�@>0	�pWx�5W����#؜"���ij�!���k�"�V$�H4�~]U���/׵��wg��H,�}��z"%�K�P~+�p�H4�pY��N�DL5�G�)��2��G�Ӗ��=�G���-����0�4�7�;e�Zݱ�jG�X�<
9ȁ3�t�g>�-e�O��.	��0��8�I6x�3�L�@c[���6:��Ueie����	�!{n�@�NA�c�1�i�p5�G� h-���*q�����L#���Z��:��:`�-@e�;yXZ�h5BR�6�W��u�K��-�z�Ɗto�#���cWF�t��I���<�D�2�SںEx�6�(�h�,*o��h]�e78�n�)G��Q3�N���E�3N5�U�t#�Ki�<���u{^Ѻ�k��Z8B��d�S��d6l����?*t׆�&e_[9�]䔏��0�4�0��3{?�t��,4]<�z��e�������)��]&�X��A���n�3���"���!_b	$��q��5ш�ӯvP��iu���c߼z$���8�^��`	�&+���7C�sf` y�w:����QL��c:Vz�Y4o��!�Yp�}��@`�$Γ����q�ɰ�1)��|D�S�0�Ē�?��V�����hX4tv����F�9��b���Z:p��D��9vz�Ъ�Z���j^9,����#uR_kNE��T^�+�����������$U��:�ߕ�������?��C��[�"����V4s���W�%,<:V-;��{5�{򰱷��{�%PD�Ns�]�,I����J�cg�)J��qk�`,�G[sT=�=��s��Ƶ�yN�^/���܀D���_S�U�j��P��P*��#��%�ƫ:��)��1M��<ei��.��{ۇ ��Z��HU����8s��@[�IU�	h�j�XFӍ^�7!@G�5�:*�����>+5(v7��&�`��� T}�c�zƱ��k=�*V:�UV^��1�<r|���[h�!u��u�j�J���݅t�[Œ��5�=u>@X��Ι���k����żK���y"�,uSm?M�58� I+�cdä�%��g���)�d�1!Ёh�#K�t��ǹ�w�02?�m��99����]�9�w
��p�.��e�b�[;K�Hk��DT��}mY~Z9���
R,���Cy�J^����o��G�F�U�����hա���pi���`��WQ_%E�6#WK��S��Jr�c[e��*_ޡ����Ufr+X-��]<:PXڭz��V���D�E�S���*6Y��Y�����A[�T�D��MmR��Bc���>Xc�~�����d���s�t��s�@�Dʰ���c��x#�(��5<�ȿJ�3���~�[��1O�] �U:�Og�5�EV���O��!o惖�[�J�[{K������R}F���5��]a�!�;G8�]�W�x �&�
a: mJ�`rG���3T�����7�z�ʆeX#7�:�;Np��8Ph���o�i|�������*�/K�\5Y�΢�Gy`^�<�%	��^'��K���
�L2�����#��s[Y�$;އڶ`G炯�1�+;Άll��� M�b�6(���d0P��̻��%�X�[�}n��nCKu��K�>��zy�-� zt�%���-�2�	�I�)tJ���o��'�L4쁺��CTu�.����:Z��_S��f8Μ�T�&�OP�ݏ؇$0���,O�� o�<�0����� ��<�(-��WCt�Ǵ�%����nM�ܗ�fG�("��Y�p� >�b�[T��>)���O(j��'�8�(mXd�7�����M�!����p(UE̠F��o�p���p�^�9<E5s�C��1�Y�Q���:
w��T�#�o�J��*I<�R�w. Ȍ_z��>*�_7Z��R�|��ҭ����-������;�����{Ծ@�{�(*(?�ܑ�K�'(�V)��W��̓mO~�sl��a6,���`~&��xoQ���Z	�R�:Qg`xR*c�_�uÉ:��/Y��!�u��$<BR���'h6!ˣ|�JQ(�9���û��pU��	�ю��ZTȍ�d.�m�mat��h+$h�:>�*~b��P�j��F}��,��H*y�.�N�y�i�֒Y��z;����җ�	qU���w{�Ze�Q�$ZU;!?�������tށc��y?ޗeu���C][�I����u>B�(zc�H�U��ֲI��c�a��j,:+wmZ����.L��+�j�{��Đ�M�Y�/�^\�B�4D>���'�@ 0j:� �Q��:*/7>>S���$���]ǒ`��E���=���I����N,��-��@|U�-�9�����q%;�Z `z̖"��=kw6wSb�z�7@�A:�${��J��e����J
_��ajk��/W^\�U��ɰL0iK�mkD�jD�=;rj�Vo�9@�m�&�{.�b�j��� �AC�k���:~\rL� 'JNU�r��j#���!�ӝH{�)�9ezA�)S�
��-h�ǭ?���/c��i(g[�����S��p�������fH���u
���ۧ���N�Jm�Ƞ]���#ڔ�hr��ˆ�����)�		"��j��¬z��N�H��)�O�����Et���?Tr���"փn?��zzl3��;���e� ��iRj�������2�m��CF��6]��O�1�	���W�k�1�7��㽆:{�WSs�%/�ҥ&����nC�?;=�kx紬JsA�M .�?�R�c?�Bo�xO����.�'����"���e�����޻e��I��G��j�x���u�����g�&�mՐ0��h��GU��NR��Ԩ�j	�ʢ�V5,�Ohv���Y��̍$�Q�&�+e�_ᜄF]�m�pDC%���i����K�d����3d@�Z�wy�	��}��� };�7�O���wK4e���Ť����@�	�''�0FC�U�e�c��|��x��S\,�f���9Jl���_P���y��E�ur��&]ʫ��{��51�D;(2?������ȧ5�z���y�A���\��O(�\w4��(�������Na@r.� Q3_����m���k�H�Zc���_�? �Jｷ����Y� A��lf��E�2���33�HXy��O�~	Q�'GHck����5L��6��ya��!$����RAv�Aaw�b�d �I�Ml���v4Q���VAη ���'���u4��B�����O�WN��|
�B�Wh�14��*zƥdڀ>�%���8�aJa��Oq�ʇDK?u��^o͟���)܎w /��a��v*�L��VQ���su�U�K5L�@J�֝g#�ӯ����Lt��2:���S[J!�h��I�ڞ��:�x�J�,�$�6�+/�4���q}A�9CeR�Y~�޺t<���F7�M��հ����oBz{6)֒P���MeX"��Z{�p��H���e��^WL�G�D=�	8/��B<��3";����!�=�E\�pC��[�"��)bH��`�эSu����ӿ����C�	O_9��;�*��(I�A���������<��E�˗j�;X��
���:�l��ޫJ�M��x�7D��̲N���:8ϛ�
W���T��v�ݕ�$i�Mw�Iʛ�
As������sU��y%�9Z܃�`.*jS��@<�}�4�M}ɗ�X��C5i�Ԝ�\ݚ�Ye%A�	�-6*�o⒬��Z,Qܱ�ؕHqi}~����?�x�qn��$5@���@ooz	�~����^*Eе��K�`k!Vrf�����.�F���gMS5%_�$�=�[��;VV��w�I��Y�6�^�rB�=#�6
�*��j1�ܵ�!k��@E�)����&�vFi!o�Gm�8~����mCD�vV�~��g.���_�|�xb�-/#���� �Of���;�b�ar݈)��#�P:�V�P�w�e�Y� ����kr0�To��p�Ș�W\+�@d�[�����iJ�e!dj��z�̥(��T-y	�w�i�!gj.~�+��T�7�Ғ%��H_Ǜ�!I�� ��k\�kM��(��|�8 �F�3���o�����\]ȵ�P�Ď
+�����a���/
����-�D?�Z9�e�����FI��/��r��Ď�K��c������OA��[���ӟʼ�:p�܃qO=���D���A�V4���]}¬`Ý���=��D"��醣�)���b�ﮁ�˿�2!����
�;#�F�N���i��=�Ĭ���5u�K��9�q�g\O�iz��.EKw5?�.m9��K��]�V�l�ϾH+L����n���w�*߉++�F]e9��Q�\T1LG�������mpZd�^�I�����s��"ٙ�m�[;����sا�\�2G�!Q�H����W��
9��h���̏�N$Gh��C�V$P7���y�&��2~��A0!
�Y͎os���I�v{��|�檁���&v�$f(��.Dt�8�⴪/5Zs��i��B�j�P���LC��?�ou[~>��^��gYr�B���]���oYn��`�31-�*��T�TS�D�f�j �=x������W� 3EL�6"wݟgZ���V�e%��e����F�1�����AJCJ��\�	=�����(�p�5���~�S��L�K�j�*��J`F�ݸ���s*^��;���{�5Y~�T���v��=���q�9��W���R�����f�N*X��ָN\�L�=��1�fʨ�l�_j�~����Y7��>�N��?s�ۤ5&�h���Q�3Od_>�������a_緫��� ��M�W ׁ����"�$s�n�\z����D��A�W�0D� ߫�||����Q.����p�hB�L>~�lEioB�rX��As���*ba�Qc�<�������ܼ�y���sQ|��Ӎvj�AK��Y*�@�P$�0J�E�a��(���x�f���d���9�[�4Ցn�7>dX�\h\ ��t\�j�]�}\���6��GhD`�죞ب�]��o��r)�ov����Z7(�X���!�C|;3l���k-w��@��CNƇ]Br9�O�.�%��t��oxBπ2��"ze�Fs����K��z���$|
SI0��Wp���S%�ʫ��R����p,��"6�2�P/���%����UF
��8��$Ү�!�q$R�m(�}ף6P����?�@��yy��c�[c��c<7$��Z��ҊAI��30�cs��/d�ӱ�V�B
$w�I�0��Bd9;;HI�K	fЇ ��q�)L�Yh�x���p�twzjt�`������c���ӰE������N'c����IQw�{���c��;�VÌ���'<nM1��
B�me�}�.'Y�od�y����։0h������iv��$������ϋBz}�X �!2@ ���A�YrK���;�9��o<��D;�>�_�^�}�Mm�C��e�����q�T�4V5��FR.�~�I2z'"O�T�rxd�2��谌ݎ����5�?Ǌ�V���L/�K*�
� - d��O-���|-����$�>��R@��1��4a[�c�*g����74�"��`��S�z��<�3wH��l�N$4"7-KK�"�,���չ�B����f� 4X��B7\�Q0��ak�kzX���E2I=hQ����l��'q�-��v��1���BqwR55���
7g�`Q��y��clk�20���=vs�6�����(dK���,ȶ�]�� ���}���
y_�E�9����G�I'Y��������yT�]�����BV�bARL����P���sZ;eg���\�\�x��%HH�U����E�Yb�H�c�"pf����T�R�S�9�]��H��o���@lQ������
��y!Bp�&8�8dm�ć�=�'O�ú@��������`{|̜��K)����͓���%�%vM$�O���D�dZ�>���rw��%�B<�fyB)�x�˧򉋴��V}���D�xZg8�����rۢYfG%�+Q[��k5	�y�C`f��F�~VS����c���U�����Rcǜ����z���� 5#ֵ����Ct��>��$����)��U��_��O�{w�w�}�hF2�d���X�N`�����C�����]~�G�E����,�e��45�m^ X�����U�G�o����#}��}��/	��>�u�^���U���w۾�$?�)�Q�Y/�1�ˤ��'˚l�
�47032o2r$1�t�>���z��L�u�&G�o��r��BH/L��/���~�r�v�}7��j	�b��-��ZGܼ��d����L3Wfr�*�5�m�i�����Mތ���+2�]�C(�~ ����� E��k�� ��͵hI��is3w�~�黪�����<��\���ؼn���^(�᣾�5��^����t�u�����.�M_}a�,���6冰���ŴUVZ��m�ZBAAc���AY)�t^���C���$�}s��q;��Lk���Ķ��D埶e�������T��i������ߕ63CPu��7�V�  ۛ+Z�\O�Ĕ�sS� �	!�Z���~6�����9|*�L��B���U[`����Vެ���2���Sk�.֢��K�(Xa��X�	#${��`o���C�@6Vb	�����R�aSb[K9��tX�KɍQ�Yh ﯾ4o#f�E�cR��y��"�����͎���n^^��U},Э�Y�F<�9X#
q��+ZRl��ņ*_�!2��$��Ԃ�uMh����v�X,Y.i���<�����$�\���_��o�T�VS���L��F6�!e�3,AJmQ�L��[ъS|R����<F�/-O��g2Q���)+K�`�u�6\��No_��1 Z����Ҍ��ՓY�yC[
t���]���ՋJ!�?��.>�I���K7��P�1�@l������b,��)+H�RN=q��E `�(����6[�����4b���e��k8��'�gz�H�y��ޞ��߉蚘�Ցӵ݂���Ɇhާi��0��я*R_�>;�A�~�EƓ�j��-#�><��v����bH锉�vu(-�Nh���4���liH,���q��3A���;�H�'o�sU*�0m�s�,�*n�sf��o0@mc��"2.�i7U=I'v���DhI�0Q��߸�M�<:UE��O^����(�R� ށ��_���U�&�@�e��U���G�I��P]�{&�#�q)�(�K�{�����bT�'���)@=�M�-��|B�\��&��:
qb�O�(�(?w�󖭪�>�����(�N��,�ɚ(?�����՚3�7`y��f��F�Y���D�u�h�Ph!��۽7�R���Y;����5BU�� ??��w���`��WL��T������>ϭA8� �0&O�V1#i��2�7���H��G7��U���(t�7tl��Xm��D`ړ�o�Y|����>%��5%���m��"m�Տ�Yp�id�eޕi7�馛���x��C<:���SC*�m��6��sB�+b$�(�ܭ(m;u�7�1���;������u�xO��z<@���Ȥ�H�(�k�K�hY��E�M�����r�d��b[�a�"I+��ݳ�7�w NNv@�޻�"ѳ�Y-�7��2穯"���6�@��%���D7�����
[�����(��1�~���~o<�*�N����o�[[L�dx�h�Bu�a/]-���F��%ɞ���� G���u�dKv�.(gJ�Yf}8a�m
�k�.��T���e&�ݐ��!E�H(y�R�C�w�G�
�.�O�r)ە��X�����
! ��v�:�X]d�y,�Gr��*Nv$����{2 ���})N�29��H�`��Ps�hf6���N�*R������ܚ��d�/d�f��A). ,QڳJ�h*�D�JQl��m�k��9�2VB]��R�ӆl����^�L���.�<��'y_�����i?QFepcB�~/	v�(���:O���#����~���?1�|��Br�b^��9wg���7�n�Y��v�&�(c�r6�Ŝ�[�� ���1�B	��R�Tżx��'�.���k;郥稹��t8�q������{�������,p3��M���c;�S�O>~��X�dL5�t�R(��clDr���Cg���)����c.��Q�����4���R�M�"��!��(rݔ4�Ԧ
R�.���uصA��m�/^�i.)��E�iFvP����^�D�<�HC�����\��ΗJ�0�$;ޘ��.�����j��|x"�������D���e=\b�+a�"@��MG��	+�'��dg1R��̶�3+h�]�5���ZM��ZF��]qi�ԂR+:O���g�����*�8KH�$@��xP_F��鼳��|K�a�!��;.�Y��.�M�Y�����Iۈ�l!���%lS|�M����!ڪ�m҅5��W"���K�?Zr7X�d�g�j�@G��/Z�����Z*�vpȕ�=�wtU7��Ω�t�
»?+,G��_��KC�-�}�h���vz�O��Pm��ЃP6���/�,���RI�1�5}�B�~{����H���!O�v��T
~�@���X�b] ��ց�a+p���tSg�(Ċ8pvf���|���#*��$�FO�iA�b��g�v)�v�$�$�J^�����>S ��=8=~TǬ�gq�3�H� ��bw5C���#5�H�`��ʡ7C����!ʲ��fFv�C3�vg�m�%c�ʠ� 
���'Z�W-`��XS O��(���K �Q����M5g��HK��.D3���-M�we�)�K(K��7b`:Z���� MD "�����,z1r��,��'[b@j��hp�hSڼ-�>�Q&y7��'��\�����ܻ�%PZ�xt#��/]�
~'���n)�n}��h�?�ZN;�)�_n���/����B1�I��=M��P`@�����W���4`�K⛶�$Tی�$�· ��}�H��$Ų'�]
"�M�_���Aw ���LS�Y������(`�Y½����O��f��]��>�0�����������lJH����_�# <x���	�D�� ��1?�ah)���s"]�q�X,��;s|�QNW�ڞ����W@�dJ]�W�����z}_����h��z�Hs,�#]�lj�����ZԨET�)1��'�]x�-1E����������L�ن���ឺE���ci��cѷ�������\X�`Y{��LH��+�aW:� K��XM�n�T�cgM��j��K1������ŵH�ݮh۵BKR2�ۉE,�'���T\mq�o�[u�.U[���J��H?�:��'=�{�����& A���Fk;����{�b�b�M>�<��)X���v٭��e��8h*��[�?���+	�L㽸��Y�(v^/�}����Mv J�����*7cN]���]��AV
*	f���7�&S.�<�A�!�������ٿ�v3���ֿ�Ü���:��`P5�bJD�@nŏ�r�x�wޏ���_�m��|L0�����FV^�m���u� ����:�n}�/ÁO+<��Z�T��d��! ��]�o��!CJ�W�%��E �ٍX	i�������k70 [-��5��0�f��U}���a 픫��V�MSȊ,�t��ZųYł��M����<��r;�e�3�%���$z��M��$c<��N�nG�e#R	��JmW*�0�;����V�ݪsX��l)a���P���K��Q�����2�x?���mL��N�3_��8��[�whw@D�����8*�<U���W26)Uj����麶�;�C=�DJ�0�bݼ!�:ehWu-/Jo,I"�P�(���[q�n3 ����b\,ЧO~�&��E��͚Z�=E�d�fv�}$�t��4�И��(��3��f�)���I��Zo���mSS�zdu�"h7�(�r�ߡq���?��,� ��}�R�k�Sm\i^cqm���
k��Ǐ�sK�U�X���n�F�� g�ޗ`���~���5��BK 1=L��Jؘ�[����J�hz*�~��I�:;�.�ߜ;	\�49�=&��{4�`{#l]ڜ��A���GS`rcL��q+�,�d�:�[�}�/Ј$��/�������Ab����P��!t+�p^
�4���P݁��2X�J��T����J�����APƂ%Z�>-2�;��.|c\l$�P�D�y�튙p)0�z���]Z�����r�9������QJw����:�(��W�c�Ib��'�B���-�tká�l|BGiݍD�`�7�"����
ܵ�Og->����Ѳ��@2��f�m[_Jv�`F��i2�9}^��8�f����'�d� ���=t���o ��9��
�}"�BTF����(.A\��su����:2����>1Y��1 6r4*g�
��d>Y�������*L@�WP�|����|��k�^Wm�8�k�Jiʺ۹��]?x�y/p��b��B0�ņJt�gM����)P��h�b3�d�@5�j�,�IWU�ӂi�Q����ު��ٳ�:{�B������])gt����e>��\w���?co'4d�Q^$�\}#D�)�o`�QO�B�eU����MD"<��N�� 6Z��Qǫ9G�]U����G6t��	�(��]�v�'��Y�-ϫ*iTd����Q��a(@n$xL����~/�v�oE�	du:���O��c������4Y��,�ya�J&#t��{�L����
����\�AϨ��2�S9'�Dhs�f{�0�i��*`�������2���F�		�⁳��-��l<�C���;;�ǈ���>ڽ�қq�m�tm�/���9\��ZK��|�0$�A3��}�
=	mS��ܩ�V����P+,���sn9I{��J�hl�� ��صP,/�_ʞl���Fe���q�d�z٘��gX�D&��v��3U!ō���֝q^&�7�<A�lY�*Ŋl�����G$�~d�����&dK�w3��������,-�!���=�� ���ཡD�f�;���B�VH,�ɻ�ό8�D��0��t�`�ۘ�2�J�\�%�D�#Pj�3���k<��a��������iDWW a7�!�\m��yΪ|/ճ�������Z�&Q��>fE1����Bx#y�
�N���>�>�XԘ}�\����� �f=e����t3���,"��J,mN�@����> �}s��I��:$eA3�T��L ��=r��B1���ws��˔� 3{Vޒ�p|}�Q�N;P���i�M��<~��j���!���)���ěb!!vw-3�����m�f�E�j�$�����g�%p��̅���������F �nҋ������фjP����,�?��b)��&Nr�w�Є��}Z4��FZ*	q���C��s�R�6+*s1�ɷ��`ne�`�����G��=d:5d���b�n����"B���]�%m��;�y��Ar��۴l�������p��:	?py<����I���ms�eI2v�&�}>H�L� �?��	�!��f%>����dJ>������-ISY��\�zlɩ������� �]%HU%|�9ȑv�f�������o~�,�z�P'��҄���X�MfiP8�������3�xaK�J!RC�?��q�^9{��Oa�A�K��Fow@Ҕ�]��>�Zu��Dto�y���[���a-r1:%���#6�b����=��娠�R�S��F���8�A�]��1���kV��k�FJ�թ��z��dRc�Si_���Yq$��-�zr�B�J�0�	J�������P��d.���|�LDPCu���ӝ1C>8�Wq�*��3���#�-��Pi���p�!����Z�ڂrK��O�����Pû
ρ��2�gU�m�e�-[��T�W��d�ϊ�B��l�_�L՛�a��գG)R�>���<���a�fp�-7;����D���ý������� ����$�c,ju� ǡ&�.�@�z��22�V�7f�=+�V�n	����a�G�&bˋ�խ!<{Ű��u���L��
1L����Hz�A�Mm�-���ewO����`v�BDDShv���:3�Rf3��?FD��yu���Xv���)���f��a���#P,dE� &q��� ��W�.�q-���0�+,��~Tb�B�i��ՊtQV�ǽ��֤Gr멎��ʐ׸��eqOr�9�=�XZ���#F���Xx3�����c������5�PEY��[��F�&o�>�����"c48:k��s�1�2�*!S�!x��y9x@a
�z&��k8X[r�`#E��<�Y��gέp�>d^c���к)*�7"�)�Mii�m�P��	�@����V)P.oݭ����3x�QC��up�\�IӜ�A��%a�O�=�����	�qES~�=(�=��?|�]���	�j����ˀdюU��[s� ��Q��^���Ҵ��mN�G�w��@z}w��H7��)Ճ�-p"m����/|eS��A���F���P�(�:���[V��f<����й6}-5�t�ރ����)�ß�늷��W����1>.X]�X��}��!���}����	�!���� �l�9LRK�ڔ!��B���z8M�U��p��?L�>�Hns	x ��'�����%�n{bdɧp/k	 ���=�󠪆��/Ź�-�X�Ss�|����<0�f�];;��*��b�ԕJzo%�j�~#!�+mZ�J�!M���@ߣ�ŏ�.�UU�>��kV���>�{��͔@vS؞��1΅%��9��bAHv�H���Xo�꺪������ݽլ9YD[�����)e�6�Vw>���W!�U�(�<��{��^��*~�[W�� ���]��Um-�S�b@�&�r�'��kV��������rjs�i�uQl���kb���u���;�f�����j�'�2:����X�/�l���0G��8Bg�s�˓ì�^��G	�3}۾� �/6U]MR�%"�]1���Z7�VK�=g�����M7�^Ldo��۟D�2�8,��Ǥ��&<CH�`�a�߷�/O-� ow���&���XKX�i��C|�v�����V1-�J*,C˅��W�>���r	�;��Àw�5��Ń��~T;[���l2��[�X�V����������*/�t�1���HoE<;z�����¼d�^�	�ܝ��������ǘ�����sf�?1�b�����k���Z7G0N��I+�cm,T�iK�F�ƝzzPe����T+߷�j��jY"ݺ��H�j�B����`���!���ٱ�x��Lv�+����L���lA�L@
��$�A�Po��i��e����Хfc6��߅�>;�W.ك:�"�-�/@۴Ƀ�{ǚ�O��{���K�AJ��R{J� ~3�����2T���f��T��D���z��O�3/�o�Zp�Y ����s� B�c�2�$QK�T:�/��(��,`�Pqz��0#C�8TV�6$���l
�0}�&+�Tf�k�/u,��7I�3�!���s�i�J���E�0�0��=EAK����&P]���p8_߆V���D3�44ΙAPU�J蠄p�{=N๨)z|w��w��̿X�H�|��I �|U�,=�	�?&��ʮ���f�ˑ�+�>�L�_�JKr��v�o�̠�C�d��30�����0"$��K$C���9���|�'�xd�CC(0c�Lfv p�?�PyW�s�!H I%�Rb�~yH��ޡC㺴	m��p|��Qt�"�j��`�$���nJ����<�.ҍ'��Ҵ�͑��M���� ճ�q��oŭ9#ȽD�~��8��:��#��i�yi��lk��0i�	���������M��	��D�t)�I�� @5�!���$��lDJ]�����)���Oǌ���
2kB�3�΢ �,Hs7�g�`�zl6�>_
B־�%�8e9�S�ަC��߹*��	�o���l���6p%F',�%�͎c���_���,㞖k#�d�l"��ţi L��7���E�s|.x���4J3�j����t�$*�];%֓�r7���owt�R���������d�?ǫ�%L���0��N�������$����m�	`�SZ�{G��-����dA�hЗq��TO,��і��i�.�gk��$Y)�ʾ�ܴ �]��Դ��|Z�k�h��%U%� �Sk�ņT�&>q�� !u2
@?C��b��q�HG���<"����*`������=�� b�b>����$t�D$���s���8���"�IճO�m��Z�i�[O��Yh-���tS��;�D�3��2M���l��_m7������.���@�KE���bRP0l��2�� �c�.Ղщ��[�.�+"Ւ���&[�`�#��ۜ�.������t��`_?T�eh����rDcq��/�3.À�-�A�	@tX"w���91/�Rm�걃o��Q�	3��q��u�D�+���c����&ƩY�=�$���~�����>���Ŗ�Y�:P�eݝDŇq ���yx�F�������Pl�a�^t$�q�{�/`mC�y�&��?��g�+p�Z���$����۠;s�vL��6%,��!r��ז$�DC�~���
�Nۜ�b�j �0�y�i|�HO-+�9�h���.�m>�<�j�\����kΘ,s7�������N�坃���d�T���<���<���8|�p�wb�P�c2���%S#�$p37��$���V��
^�ַ뿆2�Z�r��HM���Q?i/�0�5�n���5�&Yhˢ��_�Ey�鎻�U���W�N�G�1���W���D��Z�y��7\e�����D�4m>�_[p�.�+�&Q�k��q󙍠u�W�z�'d72`�ɾ`H����Y��K����~�X+uy��Ҿ���4�١O�tO\�yKh�jg�϶�pJ	�f	MaY��_D,���.!Z����hg0y&t�6n=4����%�y�ZVХޒ���%��4ck{XN�<�@�]�l^w��M��_�QE|���Ӹ�V���W+1��V#��	 &�8�#�L�̚��$f)�]�:��ȶ���u	4����8F�7V�)�X��c���fMX{�h�.*�5�W���ǟ�0-c�ᣆ:8HTRņse�ڶ�__��׻ގ���T���zs���:��b��7.�VVT��|�'(�j�#��z�9B�ė�7�D��	�{���x����o�$gL#0)E�An���M�����i�ȕK�oj���͓/i˂#�/���Mv�֘�X�N�ܒ��y�O|!���f�B�+?�R��敥��NOq8r� �W)} �M�n}`���8�����mWv���֌�hXt_ƕ�]:js���1*J'wez��t0�j�8�W��%"��^�Ӆ�g@�����lx	�����q&��њ����_�[�/��黱1�P�P:�3Jmsf�"̓����[B�����kǑS�fR�����:��[h�r�n��,>�xy��kU�0H#%����C�H�����7I�����{��$N�PM���I����� G�U�N�rX�sK��gi�;��(��\��|)'"8A$\�6��^����65��SYoϜkR6~��'j�BH4��<��^�[��0b6 �!�j3�Ri��ֳ�1�ks@B��k'�TT~I g�+[���nf,f��ų�7�m�띥;%(�.��b�m���#B��S��D�#d�T1�ҵ��9DeTVh��/IQ�n�nۨ&�BwI��&�6��k�I�_<��ì�K'GӍ��C�\��c܂�V�<�JL�:#��b>z�2�ԓ��LNݙs#�gq�x~^o���k�s".i>���*�X]f;���`P��eI,�\%�a}{��o�
U�
w���B�������N� [�N��@�|����M�ѯ5����8az��y��rOD���L�9\��.K��U��(B�Sf�e�Q�}/!�P����I��Q^kM�B� 	+R���yN�SIo�_6U%&n�?�=��8�r����=���T��TW&�k�Yj��3���[9έ+�S�GMT/��J�Z�~������g�
�L�=x@������F�=�WY�!�3�@f �J��;��օ�N3aBX/i�v �3D�L�V���)X\#z����ۧz�W"� �����%s-�+��n&�+�pb��#����f]��߅�pr�D�������iT%��Xr�`� �O-�ex!�haN��Yx��_=*� ������/9$ �V�	]�[�(R٘����k*�:V0W�H4^���j�F;P6L��i'���5�v�����C3٩�g0V�ͷ�̌�6sw���� ���{��Z�bMX$��9q���/�*ꏂ9$u�M��Y�g:�������F�-e���@��R�����#��o
�`���D�|#���@.}��gqLH������f��'2������O���-e7'r��"|0��?OW��]��0�Y"6�)f�k�������$�[�(�4�~\io%բ����m��.��V�!�5�j�>�#vL<��XP�#uEQv�J�\(�g3�f���Ҭ�5u�vR���@��[�������	Z��$P����r���wP��y9yq���#������-���>�̲�-
����p%�AA*�������`,��bPVPn����'e�R�
�X�9^)^T�g$Zp� ��T�H(� ���oB�q�7
�����`#�
��b��}��%���b-R4��ז� �?�W���qx�h)�A;�7�<
�)�Gӛ�'HR�X�t�^���/$��*�^�Tg\p�5g#�+a�Y�EK���W�^l-�΀.P)�ǀ:�E+���<g޲e'���?��öcɲZ�\�q���]�w#�&�� �T���d���N�֟E�~#�90�#���OMZm��%�{E���N)������e�T)*ю?{��n�$��G;M�?Ǖ�?�I�ޫ=���Itq�����,���"ؑ��	S��,F�N�OhLOM�P��m�dm0,W�3Uvț&�'�@5�L$o����ߘ���i��·��N��r�*X�[r���!sx���J���E����Kh<u؆�vL��M�W'lK� ��'�`�K�~��!\i$Ϸ�&���,�_����
y�X[)+я*�2I��
<��.���Eԏ0�WM�i'j��E���ato������@��K��}���8a�g�8�ӊ�$�&��6�V�'(����R�j1�e#�<��ec�P��^�=��t(J��$�Y���V����0
4V��������,�:�Vx��֙�N�H~�ޅ�6 ogɁ<���YW�d���[]s�8���%8P��W�o(�~��iG��Z�7��Q��u�_��{~�ԓ�n(;"_D�47Y�wkWU�G9�I�=1AēBx�m|�n;�>hk���&��T���it����8G��SV�}$
L�AH	+X�(H��&��q-�Nz�II��<�
���E�U�e��wO����l��{������X���>�>��p�/ݽ�*J��E98�(�T+��BB@�����	r�����mq`Wa�r�>�}��;m��!4��פ��BqXoA(���4�{��V�*�ˢ��֡׈�lol��D6��Z����Ndj�����9��^bC�^�"�zw�u���b� �+C=����S�KX�P�
C�aA���;�a��������IǆvY��=��U|_qu8�{E��Q&िy��)�op;�]���E�_�D6W�p0_;�qۄq��-Q}���^!A�r�J���N@�:�� $NLج�^.42H�ӄ^�t{���v���y�`��RR^����%�<�WHC���}Խg� � ���lfyu��g:������esN =�����T�[��a0�kgt*Vq����w��L�\��͑�F�j���FF��fF��#���1������B�y�FmqpZ�@mk�l�Ѓj��F���е,��r8ja��ǎ��D��H�D�vc�Npiw�s5`��h�>&�T�!R�>%����o���f�D��@0��3��uBs��_����(J���~��)��,�>e1 ���Չ��@z��	a8��$:rh��$2�Ľ7��ѭd�dAJrJ`�*>�W�f٢K����r�/jm ��N.���&NM���k"��n�E$��d�>685����l;�����qo�����Y�9��3^'"������"�-��@c��_*���]�N(�5�4yzb���#��V@�vQ5����Ǫ�|���*UF@b�r�^���F�����1ޒ�Wk�5�fr���Ja�i�i�˾����7cn.��d	�(����/�fO�v�.�y�ߢ���K3.a	��c�VQ֘��C��ـˌ���-�����G�];��7m`������wBW�H����i��eq��q��q��o���zS���բ�gڮ&�����fI�Gho��0z�7Mj�7��j4(�%�|0���k�Ӣ�Y�Hh�E�$�5���1 u���:!���0��ȥX�)O��N/��5�񾓇!�M�Y��3�b��;�ҷ;��l%r�˸H&E��Y�gC]&C����#��7���E�P)C�h2k��"נ0�9�>��Wf�fu�;�z��o��}SS%|��Ԥ�2]��K�ι�؉
�c�%G^"K��cE\��㵎�[��"V���z�Dq�*'���ά��k3�G��i"�v-��Y��&��$c��m�W�bpg�A	�z�3o蔜"�l����9�0��oL�5��;ڻ<0hU��#R���D["�����
�*,K�J)C~���yeu�n �ސ��e Σ�ЋI���GbLM�/�ז�#�xV{���m�o�%�q�4�����Yf,H��!=�r
TC �ᢳ���J�1�GTooBS��6)��r,/���F�����?
+�jI���EH'������|G0��5�7�'z�yG:����~L�2ѷi��+j�h)����4�Ǭ�-�5!���L|E]
A��淪FC3���m���\Õ�#�M�ˏ����ل�JKT�&?d�1DX�G���1�����J� �rF�(�F��)�%��-f�ǒ��i;M�`�۳*!���* ���8p>��o�1?�G����6|l_�]iR_Y❦cch�~�Ƨ�g�F���HgϬ�g��(�X���\�䈪d�y]�خ����
=�N���L��U��7o��I�h����'jRSi����Wd�K�*(��Ѥ�)`�ϨO�7�Ў�(F���sn�S��+�ez|;��D�ڄ�� \�m�7�� Y <&����ɻy��1���3MW�K�+ �T�|Q��s8�Zu,z�k�x������j.#&�C��7 �B�������9�{&F�2e����Yzg#غR	�V�4J6�)®Y�+L����i���}�b���A������=h����=������4�r�w\ՎJ�-���j���h���]�O~������`W��`�O+=�>�������U��/=�xT�+R�:�j��	@�P�"��3�rq��e���,��?k�$��|�&����L+"5J&�U/kl��}�3�U[-��lY;� >��F����{wLr����އh:ʁ1we��n�i5����y�/�P%P��dMr�۝�|i�>���C%���6���$ړ��q��@���ɸ�Z�8��I����`�͂L��WBGc�H�/W���'O(���.�pt8f�	ɋ#0j��4��#������������Z�1�}$���s��k
Ģᕕ���,*��q����m�Wۖ��4��:0�G5Uvl�|i;Y�S��
�Z��U��zL:�B���9�c �y�d��Wq���������g�F3�xn|B� �\�X�I��O�^�9��a_��e+���3-�����Pb�Md%/���׍>��D�K3�唹������$��D9;�f��o����9u�(��/S��N�]��/������]��J�����34cp\cg�
�)���K�BU����ɼ�*Y�&�����73���\�8,�(�a/�m�C��Q������xkٮkGu��%<�49nP�p`dm�lgf�#$\&����ä'�f�τ}8P5�����.�
u�0$]<u��!
ƺ�*�h=��=�|!@��ͺ�'V�eEf�
P�U+�"CW<= ���t�<��}{���q�������]l��]�8�<�5�������^�zm-��e���8l�p�D�ᰣ���6�n/If�w���K������&꟧�杗;��D2��@��[L�������'�E�d�0DEs8 1�?V蜁�_J�3LWxP�����h7��2?6D_%�r&�i���.�O��پu�t���Ođ":����]��~�
���^y&�i�y ��(ɝ��?=���Ӕ��Ն4<�|#�|dr|�E1�V^����C`�vE��tP�0l����,4��:G}���u9&3A3]VD�RG�Ij�������\�\�	2Vɹ���c�h����5�r�y Yf(#,B��B�R+\�G`YNZ�+ط����n)=`�TU��-Ұ6��ج(���+��T}�&u}ou�2\��!�2�XPN"B�W��L�8(��6|Q7��y\R��Nڸ�=<Y()-�����mRu������m����Rl�5dM��]�\�)���if����;�a٩tgK��<���᐀������m���t�{m@��j_�RG)j��jŪ
oN,���U�T��(���X��@�Q����B��۲�n5ш̀L�A��~�1�7*�llo�����Pi��0���Y Y-5kW\��<��K6c�c:�'�`�&�o�Av6�1l���|(:�4�􈣫��#�����XS�.9N�KBv�����,f�"��"� ��#�ŖP�����mvY� ��j���#p��pͼ�G�پ��V��&�#�;�`R���B�Y9��!�N4;�
8%�:x�B�W���c��n�	�4�N����j3�	���m��K�ßsx���t@>�*�wP�j�
����2�Ҳ���bC1�>lJS]�wԶH�N]G�N*�B���s���uɀ@\�f����2��n�f �-J�N�c2N��1��6R����N?+Z��"�q��\�yIT�g��kf0�q��[�P�ؾ�]���k\=����H�0ٗ F�M�����J������H�/(���.=�֟�-�P�d}����߱�-@e�z��;�
$㹭�"X��)��K(x��0tr#�D���^��# eU$7��&OY����J= V��pT��"��yM!6�TB�d���ԙNa��ܡ���q>K���}�X��
��B@�G�c�0�L��L>���`� /C0��.�=Y#�[��e�НB��f��L9���yWE%[a�2WƮ�8Qf�G����MQB&NɅ5��9��ǻ�����3�FC�ג�I>�yk�
��t�+Oݣ#{W����B�sIw���I��o/�w��uc�,B�9��$��ݿ\c
u͛�BR��c�9��Q���맕-�J��o�0��J�PL͙��p�zG���Ñ��Y�{�(L5"��"��2`5u�}�搋�R"�@!�Ri�=+ٴN*8nֶ��2m���A��!9�]���ê�^~	�̗�����+I���Ӛ̎GE���&���
JZ5��_$#����E��EI�9�z�cϏaI���j��{����gSC����ϵ��4��~��՟�μ[�0E���8H o���%4y6*������eȞm�T��b��,s�!�,��LT���nzQ<m5-�)GwI�:���F�:�Va��D��;�[�" �������*��썢�#G��y����J�T���%!|ޡ1�,�x�죆�V�Z�P2�l������b�	������}.@���U%mX7�Ά��dA�����{Hlh�K��$��l�GZߋ\jB����9�k̅8��AΠ��E �1��D��@�+J� �S�ME�d�]]��v��k�g}xD�'CS��;/&����~�Fߥ��Ie�eɱM�{���̓1����:��u��!{,���b#���ޥܓ���$#nͤ{O�K��\�C�����d*��R<��S*·�Z��)޻}	}�#��($�΃�#n_�g�􂍫��A�'�	�L�2=��Z.|:r���KJ������3�Z�T��=�ي��σ�����g[�2�hU���㰴�'�8]�oJ�������hK����t(6��sԈ7{k�B,&z����;��co�;S����]�vBBE�?��E�+���$V��HceRo$G����-�6,��t(r�3e��T���SݝH��w���7��_!��K��\�54��Řq�Gv�{Хe����DV� ��u�p�� �F��r��_	JI��q*���=(U1������̉İ:�����cK�\��h�����t^K��H����:��p'���i���A��7����[���T$����w\q'���)� ${\�ę'��}�&d���"��mC�a�]�J��H䯎�1��ZM	,��a���|9�  ��ՉQ�}3뱛ݿ���J>C��Q�G�AI���Q��3ò�"����]��[_��_ud� J�oU�}��kE�(��]fxB�yE
�M��7�!�ۻ�N��M����Ŝ�^�3��M:�]��k�%i����Z(T�Q�uݬ�t�h�5@�x�-�.����D%3�i*�W����<��7�~�V��C�(��H?vf����Cà���1 ���A)։3<&�ι�/V��K0�ziw�Ǣã�&/k��K��>/���W���sP8�??2#�y�֐��ѐv�fxj����!
��v t�!��=� �"�΀@y:�[����;l�xc\��¹��®���ź|i�Sl�m�n_-٠�b��_}��\It`F�U_�� ߂1u�dYy���f��ҷuH��24�َ���xOx���g�0{F���,����}eUV�F+�e+W ?S�M�� a���e��Ϋp:��&2��2��j�R<`�t�� @�$����2僇Ty9!�G�h�5�~Lxc�(f(K�DA����Td�����,h�jk�Cq��ڰ˴�Rų2�����X(we�R����g=�WϹ��fw�~��R�x�a��2|U�O0�0y7���~4��X6 ?b���B�< ��ڊ��S�f�"�O[�J�^�����Mz͢�Nqui�Z�����i$y��7@gmg������Ķ8�x�6����J����b�/"6��9@�khI�����I:�k�O�e��q�Z��ּ���k�0��BDiCٹZefi��h�2,�Q	^V�!�޾�Ax�U���v��^B�����������mGFt��H�O��e�� ё����ֿ��bV����3������ $5�kV��)��Df';�M\P}���׾.��X�ZX�> ʂ�*���̊*��u�q���
�[�?�$:w�%���X�!�2��ĕ]]V���O* �B��0�R�ҥ���hD�%�
`�9�z����&��"t5M�?Sm� S���%ڬ����
�B��'�\����w�s�֫�^s%���U��j7Ě�e�6����;�;{��%��_��)y�~9�������Ti�e�?{�ԉݬ�2�J�n�v�RZ�}e�y�/)7`���ʻ�I��{���v#��&�eO�o/HR��o���9�+W`ktT�f��D�F�U�1�.�c�2�;P
��t]��\Y�b�8%���k{�G�t���K��9{8��t\'��/��x�'�VU@��o�
�ѧ���f��$�77�rf����|~`4Hk�< q
�����$��	a��BJRl��B6���t:�o#��9� ���t� jG�������d1���z5�"ċ�K���sC	�;�}n��d���0x����J�OUL�i�>dM9�����g�n�B��]��9dw��Vn�|?��2�)�J >�<
��+�fK:2-�U�E��P��1?�%͂q7V�07I@^�I�����?�'J�[b�4$%��0M�"����M9�H��s�}aP�Fx̡�	�R3n��٦��3Xܹ$���*�3&�"��׏B������!��^�t�kH&Jk�*��})�*}�L@Ƞ�+.&kQ�)s D
pz�s���X�7oN�:�����&Pm�6w��_�J��ᜰ���;����j��X�~�NUHh�m�P���2ϘeU�凞�+>�FS,9�%h�c�9�j�C�[���gꊫ&��CȢv�ԗ��MC8���]�0bE��n�i�U�������J����l�E,�Y��I�X%a�u������bsЁ�s�:�=��re��}�4.:A�(х��)�~䒞��.��m����-dO��PgI�G�:B�uq�e����c+���*�Vr2 NI�L��Oj/�wH��e��uB�L������y_s2V��t��	d��_�%A���F�cW���Xc�͕�16��5&G6���Zu��xیO}�	�ԎL�|��6L�b�9�5LWNҠ�7���,ɋd��sy��^�C�5��<�Ħr�I9\��~���M-Ę`>�ng�KH�0�'���Y,�z�>��,^Z�S�����Ƞ��f���
h_�(����s����&*6Z٫���_l��%�C:�l &$����tx�QN�M�S��e�B1��˶x����bE�������*jxg�봡%$�m� xmƞ9��h�n&�X���Mp�&t�ܩ*Kt�����x��s�/1Q�_8����U����}ad�:-�<�6�BK��W��A�@���~�i*Х�2�)��m'�Ixs�ٯ/V��]�!�gŝh�p55m)iP*`&�xvl�Rޯ?��c�)zfR�l�d��#�)��E\~�w�u���ӿ7Y�r���>�D&�ˉ�=����U�ǫw�>�������[L�Ρ|]�ʅ���#�G;eǬ��Ka��<���
3�� d���ܗQ���4�w��J��8\;�H�<Ðs���;�|}�.,-b�ⵦ�z
��~�9�����%����7�tˣw0햆������A�}��%]#�n᚛��"���g4��x|���9��-R���%�şȆY7�)7F������ǣ�<~�Lo1e�m�_�����]��)kX��V9�	�Ӷ�=W.����#�/ل�JY���M�:��I3BfI;v�c�H�q�L@����)A�h����T�;��%�_H�t`c���0f%��gpbߋaR��j:�Wǋ4U����#<YԅKe�?v@̞H5��q;�ş7�<d��ޏ�%
������w���%i!z��ǜ'&�b�U���X @Z˚ic"J�+;�-^hFA��zW�J��$�C-�diG)���ꋀ�7���1b�	Yi,��o�RZ��u�	�xS����1�r�9.6�]MADڂ,�t�����!��S�G���m��|.�?�m"�l���a�ȝhA�x�~L���wxp�$Ȉ�%�*۬ÿ��m�{t�P���5|�}˓�����H.I����J�{a;�
�r8�DJ�4K�VE0�Xl���E��3���� :Ԛ�;T����/�]/Ew�a�vQ���m�e1'�l_(�\�`�j�/�������	��>y��a��8��|�i҂��qv�?.�x1GkJ�/�ˠ|N򑟘?E#��0�6�QN7+����FI h{��g��hV�n�J;o&f�??��7 ���09	a�(!ن��_s�jN�}V��8j�����
�+&5�k�b��ۆ�AJyP���.�#?E�?\�x�崥��\�ڵ�-�q?/�}x��(�Pi�>�umwcx���]�D|d� u�b'Bs	R׋,�:G=�y�:n� }���UU�~FM�a>�X�������N�(T�/G���ARL��-��q	��)������wb��CA\�F��]�Ų��L�_��'A��&�u4���/Z�z��j���c�,S�z�'���م�U�2����e�TH�'oDN�
���*�w�ģDʯ��;3�?��H��b>튘4��R�O\�����������X���`��^S�`�� sAč�l�w��rnI��m!�\c(�[y���{:*��~����� m�_ܞ{\����M����R�ښa�u�U�=����^A��U�͝�Qǧ)O�,%W��Lld^�+�D'K���؝S;8U�	v��~��E�C,�4���9��1x���Y�#,�B�@��R:I���%tK���g��/,c�23d*�p����K��lB�LOí_\���~�֣���f��|,��	��,e�
_~[�q��(�j�瞬��_�F��e$�D��;��\A���B<�����6��3���-�Շ��S�t�=�`b�ԡ�}t���C��I�P���ϩ���o�^�Ub4q�l-�,Pz|�`���B���T�TN%��Ǳӈ|��4<[��RZ@�� ��g�AA�G�c�Ư>�g����\zDQ�&�!B�H�!.g�#��(�	�cW���k��hՆ���Vu�lV��<��]��0���؁��uh��.PV� ��{'����s�qEƉ�Z�!b�3����)i�?U��;r�W�V	pW�Q�Kd��B@���?�tw��Y@�3F�[���Ք�֣يZ�q�_�]�7���>���v|��`��S�\����{:Bi�� p&&|=�)^�8p>;�A��I�D�+���w��i���2*�^�V �:��P�<��7��uz�9�>.^��7�b�`�s

-��/��M��ܷm s��½�O���(,u����l{����!��`�0O"��mQ͹Y�uuzUN��E+��Z!����AZA?�L��b~�i�{����YC�	c��X߸���$Ŝ%�Q���؄��!u� �ob�}�FRH���W=m��&C驹NB��b��r����hw�]�M��A~n">������:>My�cvlE�F��x�:A,�p�$L�K�v�ui��J�;c!z`$f����{6x�*�f6������<�O�S>����Y�����*z&��$��K���I<K�"��N��y��˶��`����G�y�r�3;���_-�ݨ�]$�hz�9W��NP�fe�0K�@6��ߍ�X*U��)z|2�w[C�)��~�$.0���铽�߀��\1�_��_��������1W�@J[�wSN���/5m/倽2�Y�i��u���l�w�e��M�KӸ�pN��t��?���A8\3�.�8�d}��g��y8�)����>�<i�{K��j�v��@�����z�G&E@1�EL�A��uǕf��'�C�A �����u�*�_��1*�e$�������3"�*8��kb��h��` �QCO�
𻕀
���p�����^.m���'#Z1�����Md�We�U�W��Xʍ����l|��J��G������A�*NlbC%ׅ���6���)Qz��ga��>�7M�궞3v�R/�3�淂�yxt7}��z
 �{��������"�6�M`,��pe����勌�e�끏���Pi)��y+��a	���i!�� ҡ��a��a������}b��x.n�ʖ���ixG���8�@�ݟ
�%SI���d��j( B㻦u�td����hb�lIxp�=U!�OS�GO�x�L=�����A�+���!1#UE�z��%�'jpIQUvSg������s�U̜�p$z{��#E�E�?���[yE�mMBz�'��YY�ĩ��O"D�=)y٣���8�n� ������cA?N�}��8���8zrG�sLu�S�W�G����wf/��n���cN��M'�u��%x�ng73 �P���9�<!-�TD�2���ޟ=\���H��%FfM�$�a]-��U.|�}{��s��BOwm��*�?n�D�,ݮ�����'*��;Ȃ���r[��w�=Z�M��d�H4�1m$��#/�-��_qڋ����8���p���0����/C�+_$�����C��3�uO��@�5*w�C`9,|
�R�5�1J ���3^=A��1�|�#BBM�����[�E݇��'8��hW������ɘ*-,����&�N�K�I���f*� � �6J��d�����1v�8��v[}�Ť<68���ˬF�e���	5,<0���$x�~a���̤��@i��q���6�^�B��/�z``iwO��i�|���6ڜ� ��i�,!�ڤ�ܩ|��+1�:�/\A��ˑ��a)��G^���ys?z���*��^�_�-x��-i���F�$�D$i۹��t��rH~<��I�F�M�ݜSfD�������m<��,U�����~���Ү^����d�%:��
�Q�qGX9x��@�_Q҆�Pj C�'1Y�K��%�&����2L�r��"��G$�狃�ރ�`�'ZӋ�w>����#���/9`OnN.���벬g�6��
�3> ~����Fbj�51|v�	y�,�B�(7�*24S!3/�����6dy��04�T�J��ODP�����U���x�I�a�M�4����dd��7�����(��L�"����q+_�Wt���ܐϰd�#ò峲w�0+E8��6�tP�3�k|�����H^���}���H׀��b/�%1�uDʗW�3ȑCNGJ��$A~ic5�N���A��Lz�B�9��7��I�֖u@ZW%h {$ �<�[�Ƴuv�_<�N��/@H��ŜB� Iu��1 �+�Z������UpV�4j�Fţ��D�/O�"g�/�!*-�]��帬�؇�;�n�po̡�P�"W��݃n}�|�VIU��	%}��ǥ���oxNL�E�^/�>�3k�O��c6r�z�㜨�Iz��ũI�_��D���	�Nm�����a�:��f�P�Hl��V� �t �o�m��u��;�B�$k�)����=;��*5���~1�$n%E���~�H�� �EO����g�Z�~�̣�-BSvo�nI>ĵ2>�;aE@���S	:')r�nE�R-H(��'ʬ�s@�\Lz����\Z�{٨kU�A�
g����2��i�?���Q�8"w�!1KxW6?2���ܾ����b2⯞G��V��&�P�5���Z�ū�$����G!	8XykV-��:~� 9~.��_5K�|�m BDT�$j�3ً�%,
6����7T���A���0�R�/ ]�P'͕�?�� *Q�P=Gd:V)X�=мW��)�W2a���إ�o�]i J���Z�DzR�Rt�Xlܪ5�L�'"�YG�LT��b��b]�ѿ�� S�ݿ�C��!�?��/i/�z��c0�j���uL��?���J�w�,̈́��g�Z8��;37�.I�v䲰x 2�܁�ƊX�ݧr�3=l�
�p��s/���㕷ze���D�	]����*7�sQg�����'��s]��3�Oa IO����6o-�aA@�߾V!��P�<�kb�b?�;�&M� �jX��R=�}�KRT��
:gg����[���)�Po��sAN>ą��=#�!��I*�KYƔØ˟��C�/�V�p��t{�y�7AާX`7,�<��E��d���:��e�i��2�"R-_�B�mrj�`|�p�S�W�<hn��B��0�}��w�����ֆ�ވ���Åy$?���.��Ho��I�5D�n ��Y���S,OS�^�KS�W�o��}˃ݵ�V��!sF�"�K`��S�E���2������L�-�V�F�ۑ-�"� |����T� �P�N7ó�1fgD1�+�}���Y
G�Z�*{j����>�-����:d��+咱�e�uC�,��.��N�9�) ��W��jV\Cn�r����?U��{�.�K�������!�P�&��N�X�w���H�@��,ЛI %���u�7 �9�o�k�
����'D)}r;[evO�?o���Jn�s\�m@Qۭ��rLx
����q�<?�vYku��t; {�������m�J �%�ڌ3c����y�VEj%>>���V�C����$�F�%d�N����dm���Bm�WǱ��n����Z�Z�bQ}��+~԰�Z��'�Iw�f'�Q���#)���"L���ʦP�<|�*b*��P\}�y_[F;)3{�]E]�ᑇǣ����h��r!����aNY�7�a.���}5���/�d����U�*�-A��l��������%�/���H�Ȍ�=bP}P�7j<���,{Z����NԤ�x���0��<��#�c�(w��xd�%���o�YI�E�]��r��;q����ӧ�[b^�����m=��Z8\��9�:��z�3���'T�����Q�lW2CT�`�����QBKI`s)I
H��մj"1˶�S�1�xϓRI�D� [�Yf�+�S���c��H�" ��E���rU�^&��:ܣs���g4�%��������A�Φ�����\�Yvn8F�M��yՠjOF�F��i~�m��?(�.*FMO�<����}��~-��v�0:��{��AX��"��/���/99�֠��.��ҿ�r���vB��!|_i}X��L0���/J/ԍ�hf���os� �V�6�$n���F�J��H���l.�$t&j���W�)
������.���/�c�ٲ�h� �
���dkt�O��J1>��ذ�䖼���Q_Fb���hj�T�9��LEN�N�i�qd����Zu�15%6���D���?�PU�x����[����:|�����5��ݽ�쪌d��dn��
��F�ӡ!�3+���mo6k\##_�j�`�!x�ϡ�&�X��]�6f.�;I`�˜x�ıe8u�#���b O���r	����c�F��o�^[�X��}���nm{���9����9��*(��m6U�#�p�F���D�H�_DP	��O!�-�uUb��&�8���!��5
U%so?�B�����&�W�1`:���_Q�}k/�7�6(��b'��*��Rv�$X�~� 8������W�1{Gg�y��$CH��̶�~9�N��I�[��g�*G_ܛ���@bL���͠�!,v����ɍ� �o	��/�	xQ��i�R+�Y^��%�og=��Y��%WѿL��_Σ� X{�߇kr��s�W��f!�(=9Վ�֛;�|���v�t�R9���p��AovO�s�7q_���"�{��1~��{����p�W
��7������-�T~�l��F�<�ф�з��8�����\X��`�/z�ۣ�
��x��<���P��M�ؓ,���B�#'����e�f�h��I�Č�9`���e��?��#7���!
���ȑ��ֹ�˙�M� pZߙ�#੬�?=�7	�G�O�ـU�����FK�,Ճ����߸�m���Y4��o���ZǶB^��̲k��`5-C_���������.;i4�8D絜�6#޾X3���|�c�9{[=4�\8N[E-�x����*�<��6An	pCî��4.�n���`}��E���1�Q_�x�9�j\�إ�0��p��^��-K��:���<*g�x��X���ܯGEǴeA�2~��e'����=J�E�$�@�^�
����Y�ž�e(E��U��ʪɡ&x7s;ɴ�8!c|�ƖK�l���h���Ѣ���ymu���^Bg��!$tzN����{������͂8<r������2o�4V�f����E�r�� 8٘t,���^'�b��[TΫ6O���,E���y?��g�p�E����?�K6.�{$"B-V���e��sl5���b�\��$��wB�o��8�����Q붕Bp{��YW)��F��3� �X(�.YW����~47:ou�/iN(}|�ъ��M
N�,��m� ���f�jU��m��?x��uŵ�d�ۍ�2�!Am89^����~^�M߉9�<H�������ReS�˚��!+.M`�x�/�:��Z	]��ph�)oj��8Q��'\ڎ��Q)G}�p-Q��V�.��i�^���=�&�ɖ+b��X��>!א���9�H�W̗����i��K;�y�枊�Z]���?�������2veS�a�*���\Za�I��t-�}o�@j�m3�je5�O{?\{=�T�#vمT���/�߉6B��=�T�'�����|�V��B�(��q�eИccZ�g���s`��ƲV��ˌ�ӕ��C��92ە�pK<��]�/Ҿ������Dŋ�l���6�=�f�#g�*#�]��?d��Y�I�#� i��?��b��+&��%���"(s�$�9|N�~���-#LW��Mz���d����Z������r�k	|� 5�:����0�2�R,��C��rfۼJ�O�)�M���r�I���|��)���-�Ibd���tY`�bĪ��)�ў �R?�6z�|V�Sb�l�S	�G�g������<�d@�XK�Ѩ���hB& m��A�<\�P����5'1����D ��ND����v2JqՔZ �-���
��O���1Y{��	��7��ҩ������w�{��|��E�t���;�U!��@�I� 2�/E9�1��c�~v�T�v�q�y	/�!L���z��w�t����v[�/���E��:w�O�\8Y��}�K�b�A�'�_�@%q�g�Јf)����M7�}/T&v֠ZI��;�:���֖ח��G#v�����q{�$"��	��L�����%0��3�& q�V�{/v!,�R�42>0�/����6Y�֭*FF�q��r���>�Ǽ�fLZJb[ڌ	�o�7ַ��1��\��J�����&�0WP��Z���.�L�S�k6X�,�YG�~K��X���U%�����2��mm��>6����C����w-0mtoO����/�s���o��<^�m �����e4���P'A� i�v��}�`}�R���ւ���Aʚ`)]3��Y6�Bm�C�8�;7��s��2���`��}޷U��Q4����I,O{�-/�����;֮����7�:�5� K�M�/��|L��� `��sd�=�BP��P^�L�����_����u#�[�,M��=�`�4�w���d���8���*����n����*R[�1:+.?Y#��7�IK�����/Z4M��
ax%3����<��Ǿ�~��ߪ$���hD�3��i�����a�w=��ǲ��c��X1��#���URJs ���2��|���K��(1f8q�wC�}��s��]�|�a�����<Fb����wRR���1�qw��vߣe��]3o�0���$&�֮C�W߶�)��V�پ������D�O�*�=|z�&��|8��šp���w��ˢ��q�@=K@Ѕ�5��o�۬D��l���O�G���C�m��~ N\H�w��q���F�*��Xp��n3�pv_�mU��v,tCȴDS�?]y�X�-/��i��8��A��:M�n;�C��k��=�����.���z���饿m�c0�b�htsF�������	��:xzҿ������&y���U�\�\�G�w�'�w�_�}~����������F�HiB�