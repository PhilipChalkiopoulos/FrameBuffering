��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾��"o�x'����ھqp��鱃3Ԉ�+���S��xQx����C�#^1��k���d�P�K}��Y:�}�ۏȑ��mt��5B�qň�w��I�H����+��1�g��x�d�q�+�+m��~�����\RJ��)H]ax�K�D�36F�����R,���/Y�����O��+f�6��z�<��Q6LڄU�:���:��-����*%n�8��B)�W3g�KEx>��m����@��w7�s�yrO>�&Y�`/��q�D�V�	#Qd-���Ja�w��gR�'(�ͦ������y��@�v?�~�)�`DP�6��	ӛ�s�hSK�y��5�c�zy,�:��7��eF�#�`x��Ưӊ .k��ɗ�� ���-�+:E�>|4�]�+��Ë�ņ�K$oj�Ra'��r���`w�d�㲏UĒs�6q!��[:3i�q��0���
�&6O��&��볁�}|�c���B���ma<M��l�Ԃ8~�������0����n �_�P��~�E�	�KOZ�4�V�L3�c�M1w@v�7�(��`�Hۮ}���#[�%QVd�ת'p�!omRT�(��y���w�wρz�?7=�=ϔ���m:�줼�'���~�C���"S�ɼ7b������-��0b�T]$]\Cl��]���0�q�̝�*�EH�:rR����~�2J{QF��T�O��y�w��G촱O}�[�g��;���UZ���2�ĝjX���y���}�}H��R��5>�1�\^]��~��Z�x�eTc(��(z2�p� 3$8�򌞉i��#�Ӌ�]�i�(�FKT >����M�=+�wI�@Rt6�l^0w�:��Z?q��E��p��gQ1�9_!�QLޣ��=�t.q�!�P����s^����,
�~9��19��˯�:RMx�8\b��r���y��4Vy���þ��� ���܀5�r���&��g��:�l,e�+�� ǷR2�2���y�D�L��C:�"�!>R}�2aoW]6L��(��t�����m�lƾ�+�<�4a��D�`�R3��,ΞI��q�ts�U�5���G	.�uF�#NcN�|��ut7�F�+ҟ�����Y4*���]�j��dM����j!;��b�zP�&gz>�)E����-��
.�i�!�t^���:�����"�o��L� >`I�i�i�eS<��Z[l��_xYr��J�f~�{J燢+m��Infװ�����d��ޒ���Ux���L ��C��YL�GJ��t�٣��xsՈ�:Gv�I�͛�162���������«�F
���Ǵ����G�d�?%6z�h|����=
��V]��Ea�%,�tW��L����Cb�l��#(D#�H��@PM����Ǟt߫��X�G�g5�>ڨ��*M��_����h;�#�,�8��K,�����K��uc^��G��@C����v�'�_�L�Y�{{m��#^;\V?҄�1f��U���Bb�y�<bgxl?u׷�\�'i�D��P.�\��V!R�	=xVL��U��(*荂�H�'�#/`�<��!��������U��\ ��n�� L��cG��3>�� g�J&6h�?l�o�.���'��2�ԏ�f�p���a/ܠu��b��)��G�`J�ש�ث�ԫa%
D��'�D/�ǥՓQ�R����ʔ���B�:�X�X��퐝�x��AX��q����d�����g("�Ap�J��6�H���'湍^��l�Tǈpa���w+%���t ��L��s��dx"@��0�*���'Y�����({B�8Y~88�M+�A���%����!W��l�8U����_�5g��H��J � �њ���.O4%�z����G���p��C?f�rG��~�r����ۚ��V�}����!7�,O�t����U1_c�1\�����"����q��0|E�A�[�'�,]H���v1_t1?UC���,���G%�����_g0&|��{!�����8{��`���;���uyU�yi��C�{eC7͑) }����_� ��D]F��|2R���u՛�P"@�2���k�W�L��B����"��j������U�2a)����XR��\�s>�j8fP�x~c�md ��#��8}{Vaiư3'ߪ�.�*O4�Z>w*-�>�����y�4���849T\�e���k�≗U+� ş���$�Ƹ�"k����J]����F��~�)���;g�����wV9u���U��,Z4��W��!�mMF�X����6���J���LxS�� ��L�S�sv�I��
��$�N��y�1������X&�����`�9����)a���]g�&6̉m����l��:��<�6�p��c������g||J���"[���1���k"��5���T�+.5HL��"�р�n㶿�o�Lz��=m9������M��U�됓��䄸X��xkKM2�l�*7f��/�9���	�aٓ�[����r�(�!
���a��yhd�� +@F�������T�4G����}-Z���]h�g��[k�ɛ�I���/��p-�A����;�L�4�>	�dM8��0�An��8�{��4�+����7@�~c&)W���n+�TY��`�����M�S����v-��#ߦ|V��.^�mI���������v��ŋ�wӤC/S�[m\�<�{eS�g���T��:'[�5L��J���q��{��
�3�a&��)(G^:Y8����V�M^� ��Mݩ'i����ZN5�RDׂ��+��hV�!��}�jL�q{,���lҪC�5����l���#��1����Q�j'�#R�b\�6.�u��y�C	`��9h�R�tY�I� ;Ė ��4*��;j%pI�\T�L�P?�3��gU#���zr����g��S]�&P�O�'�T���:0����3���ˎ
��� p8�'�8��0X��Y����$�.�f��Y@�5w�/S�oQ
�T�4��b*pϗs7nu�R�~��
��U�]DA3�ݭ�4�U�m9����셔D��b愤���$�,�w�%�'l�T��Xj��E���0l�&�����Yx�����Z]�ы�)����C_[���d�&��Q��E��Ȃ�O�P*+ޱ�ۇ��s�+Y��{��
�F����&a���wM��r	�z�5�m7���u�Tm�b�o��)T�ڬD%˛k8}�=b��n�8�)����]�_XV���.|�?y˰~��y�H����.�f�����|�䎲 ��ޕ�"Ҝ�>y/q��8~�W3%�B���F#R=ۏb�X��[�`��5���q��<<�Ȋ�&ǁ+�BR�!%���1���a-Ѿ�uf��I����Y�痟Τ���wf�}Y�~8L�E�̠_rـg�q��G��B3�x���Bm��6s'GV;{ u�83;�2"�ߦ�u���ؙӯ-Y�,���bN�LO�[��+���l� ��0�&�7��r�Y���.��	���-+�۟�y���%��%��d���R)���69?�˭M(������;�}�RB;$���C���l�5�'0ee �q�Iyp�ۄ�&R�^����O���[,�i�lDه�K��[C��"V�o���\�aG��įK&m5�,�I���w	\gCp.� �c�쒰r���@_bwgz��,П� �(��vQ�~a��M�L§�i:�L&���D� �.��D���.�b��ո��M�zm�(���UN�h�>���<8m���f�{SxB�����>'��.fv�����^8�[)k̩�4X�i�{����&��K����)����͘�^6\ҙ�m��O2�+������'�xөD/�dp;�xv:Dг�g��k�٢��m�W#!$*6������W�A�:����}5�T�L�2z��:��9�3��u�uѮ��`�r"1�Z�5���	 
����6e�3��cC�9���/�U�*�ww��l��-i�V��y+���p;�eMY֒���x@�l�
�f=P��� ���hBlb�*�:n� ��N��#�v����I
�i`'ӸH������pb��G��~��P�%tp`?j��!����kX[j�t�Ύ�M��Eq���}���t�k 1��2��Z���S (������c����(���E���]��d'%�1�N��肉~rCuS�AF�}&���������m��Ff��b.���}阗��-㷙�ܑ�q�'�#F�)CHkr���hЖ�{�h� :?,��֩egY~�kLL�,X���7��N��j�8 ����=A��AA�[?���]k�������u�Gy���t��B��`m8��И5�����ЇAK�����W�F�1.@�	������
B��!Ԕ)�s�XĔ&@���|��3�s��0����AU�I�:#�|.x����C��p����[ZEᡐ�q���)*�©��i=�7���>�?|s����h셡T�L���&�����7�C��X�¬
�7T
�\�q�&��u��!�^�hF�V��64!���O%L�e�@7w�)!��v!���o��������tRZh�TĐ�A��.��Dl����o�� �w�B�R��ڧM�5��,h��X5�o2���6Kl��;fk#��1�{?�i���uDna��	7�*�#��/�������Ad��X�_�F^��v`�3u����)�����9er�!|��Wb���>����5�4��j*~�e��;!cT�.)#��8��?�`�s�k��d$e?,�ʶ*��@֐�%�`�w��2h+�KS�@u�{���P�ٚ]�x��L�K"n�h�������t8��9i��|����/'uǧ�����-�O�D�U$nw��oA����"�K��}5�����q��7�K�{J�ʨ|�J����S���MZ�DB�(�a���~c?�cVW�^켻}`ݻ�c�j6 T�6��.rV�v��?�8�g���-g��d<���ص�lz���u��l����1!e�9��i�A��47W��Via;6�7Nf�|, |��5��_�"�����Hh��j��-��{���RQ����.�Hb�=���֜!��m��WKU���9��b�,8��S{���Շ�"�,�JU�Dl\HHn/p|��1�^���/<�B� Yr5�7X=t?*��o�ޣ� S<�;ch$�5�0N������G���
[�֌����G(1Q�I#�� Cj �o���٧�42�P�)���kCnci���F`*@�B�l\�������̗�J�����v&§e�|,�.wb��R��ÓZQ�^Uϸ3Ԕ�YC�0������S�NB����4ѧl�������+hW��%�snC�hȏ���R�x,F��jg��K�����_jH��]K�����}�m�b�;�]�=�#�చ���&_���(Yh�qy�d��¢��
_Զ����cʗ���?G`&&xv���p���XuLo^����N�;��jb�H8��R�u�P��M�`v����&A�Թ���(;��I6�~�n�2�AS��r���?�'ԨmP�qh�Jub�n���c%M��ǳ3���ַѸ�i�+T��L��ڵ-.u"�[��������oXm;���m{<Y�\v�*�-��@���+�Zƙ!Z��7O��ޅ�DOU�78�+`ta�ҟO�m��o������˲�d%�"g�t���Z(��YT�@Y&R3E`��'��:lf�	
:�܆I �u��Ϫ�*�06��X���c��?�@��b�h ���¸5�J�t��d��بC\�v���1;6�Zmws��"Q�EZ*���?Bn�?0!.�${��;;J��Z(��B^ �oz��f�ͽb5:�߭s��P'�e����O�.�c�hkW4٧'�NSu=]7��d"�,4�*0ğ�r8�qn5�5G1��y�\�w��G�F���V�mpԖ��]�229��iY�]*�F޲	B� n���P#�A� ʄT닙�y�&6��1��W�.R;��v���B�%��n,��� �/g�mcɜ�dҒ]MZ�`�G�n|�R�V�;W�٤-�ʕ[K��}�8_�G��[���g4����������o�N*�TVr0�)K�fg����ˆ/�w�������O�R����+BW�o�j;c�Ex����	S�LvNa��*�y�g��{��'E@�sf�u��I�]K�o��vd�Q%-��H�T�R�]Qc�ɧʞ�+�Ԍ	�[�8�kz^��C\JZ�R��b� n~���ѫ;Q���������1#����#"�eNz��RSV�@�E餈V+~�!���+�HL�D��=�>��?bUkGl��	�q'�VFgY;���|���ts|^U�8-��IjH�r�Ki��(]M�Y��_����8z(�N!�ۣ�����)��1KD>c�T?��t�?p֭/�rEu�n!?r�*I��)roץE�gg�,P�H�������
k�������B�?}&��YZAl����H���A��㗩��-���ENR��`���Ʀ��^�
ٸL]u����`�]ކe�M[�͒>ߎ�O�j�3[�^[+��M4'�an4;�_'#�`R2R.�d���/qo�����iDv$Tv�_e�(��Gq*Wq���G��fv�3'�$��ǀ�=nr�t� a@g��D���a_\p����Q���r�>��˖��-��#Pr���� ��e�qO]���S��]��׼#��\���;�Cs䋈��S#���Z��LҞ��c�܏(豳hIpLr��7;�gn����s�Wk��R��N�A]�)���3�:6^��-���p�k���"���d�ܞb�>I��>2�.aT[�5����"s ��QO4U
K�!��d�0��7d�fI3�w�^P�yW��O���E߿y<�;��56����w54^�%��O:th�Z��*2p�]��[��'y'B���=�)��峼TS@xz0.�0�:��:�)�J���c��{p�⶚�?aI"�UV���}�	5�o^4��yZ;��$����p��0���?�S,�KI��w%�1��)c�ۈQZ��������⳪%.Nx�����Xw��бvK0@ot�� |C9k��X�"�ޜ�\X*�����c�����\@9dv�����3S��Y.3gTu\�|�E=;���
��G��n[���\�Q�S�B�mλX�Q�M�xp���/�;�-@'���y�ٸ�2�S�)�*���Ӣ�lGk��^h8�)���^%ڂ��`���m��i��ܹ��3tp�jߋ�b='3K*M�q����q� �g�ɨ�!f����!}Y�;�iള!g�!#Ma�T��ne
�!����<L%ǒA)8�����DA��C�ꆠ:���9�˓.qê�5Iv� ��m�in�A���m��wmM9���Q�1�)�$Hu�[���M�u��~My�J3gy�R7O�$Z=x�걸t���6��Y����01���7�����/�����������wM2�*`�VC<����2�&��|���_< ˷J_�WZ;�������du�j�a���Zc����s{_C���y�d�]��Q�����x�ԼwA�no��{mT9���l��0�3�	8��g:oG��蕶TB��(�Dd{��͞�C��%����7A�4X��}
��\u2�{�J_n�¤l{YT: �%�I���mDjԪAfAT��rWø+֖�Hx����)�{�i�P8�����3X�	s��H��k��ǰ�������$۳�Ƚ�R>2�Ձ�u��N������ƃ�<2���r{�5De�=3�����>��2q�:L�ϩ�+�NoK�4b�?*���V� P����-���$R�m�Z*�O�t�iɏ��/t��S�Gňv>�T4��6p�g$3�'ZM�f��88��~��q��~<�<�>[V�@*�=+�c�N�1Ҳr�Yeߣʏ��$�Þ5!�:D߻{���=�W˖�[�1jO�s�I�G.G�T���ۚEo�ÿ `�T3��K!����g��Z�u�n�Ţ/�/@�"l����S�CL)�?/�XZ�F�K����ϫ�f*Bw�Zv��$%�*��/�`0��K �5��9IP���9�� �Ë�q�~�����:ͧ�eY�+��/0�F�d���sH�Q�˯=O�i����ʞ��- kp5qz��H��mA�������GPn����b���W�M�١��'�����U��1	U.�I0��O�3j�\�u~h�������` @	� z�6M���7����n�����8���h����(O����c���^ҹ��5����qH���e���P��k*ǈ�r/��ΰ��S���";����H+juMx�'��E��� ��ޮ"P�۔��,�-��S��;��i�8G��+w1 �}��^I���p�D�T�zrY��XH��K�%_��|�oj ��[4��|����
;%�uIu\�\���.��z؀ᐋ m���^�\� 0?~�!Xl�����|���Ir߯��uwP��'�`Q�ĲNpȋ��񏮵��))�����[%�6!Y����JذR|����k����;������Ș��B�G~`��
���w3��7Ҁ�8��pG�����r&�q����FEn�Z�Fֽd�z���Oe0���]���3�(1����5S�
@�Y�#�~�~3�XP�&L��k5C��v�Iz!��؆�g�+~`W��pmr�]�Ү4(�x�&��򋆄O�(|\}\m��n���j��w_}l:eG�r�z�)�����
��D���+����~4U�3\�C���3�ɻ�nb����i���7I�,8�]�J?�H���k��� a�^NuzAz��$ �����g���KK����70Z�b��6��ѯ�1d��� ��X�Q,���LjӨ��׉�FxJ%�/�SpF���z�V�{=7*��d��Y���׏����DЪH��4�3:�0�sm��_!Əɥ�Ӽ��bͭϫ��(�^��}jn�rN��۠�,
��h@g-��#h����L���W�L��	f(+"U�7����-	I
ӕQ8E貖���Q]W��Ȁx�:8��c�T�hY��E
=z�<�f�>�j��n�"eb�x��/��٣�*�1s�*J4+��x�3��B�
Y{ٮ�������؝��������E�F�^��Heщ5�nx�8h_�gf�C��s1��~ T[��T�hݗw�+���`��C���T<����k�V]�m ���$tߍg迎J*���z��dN̑��La
�W>OƑ)�r@̈�|�r}���({�cOjqB��� �G��MB�B���R�u��*��"ׯ+�G�ǜ���r��wob���&�'��0�FQ�A�q1c{�JHJ(+d�U�x�+!��g�P�̓��	٢�*V�����=�Yab�u�&��6
#;+e�l�����)��ҹ�?�(�N^߄m?Z�$zl���D.�h@c!��wv����bG~���3�o�t��~u�+d��/�C��`�ܻ\*���!��CY
�\���\M�f=T㬓�[ ��/$w���?\f���äQO���2"�����Z��.���OL��f*V�I����o�e}�ִ�=�O�����-r�בä\����lG&�u����,2WcWF=�������~}2����8t��g?|~-����BK��H�3T�F�͊�}D_`|�
��m�[�'A=�$�"r�95Z��+���(�\Vx�k+(�&���~��	ƃ�iBخ#X�"M�J�8��6D�fp`�Rt�Ow�G�K;��/Xt�����3\;�3'�T��oq��������\4
�*�A~�t�M
�M10�s�c�� ��[9�n"�l��%|��<�χ�
���zT/��G�j^Ʃ[s����5��B�c���^��Y����eɿ.�*�B�=g��Q���G6qΉ�/���.��n����/��S��U��52$֯�-����8����e�i��<���ल������w3�bbV8ˀ#8��C�
�����#+O�YR��c ���xhTcÒUF��F����oA�vD��)f#��THjj)����t��M��a7�y�ժ�t�R��z�$Z9L�٠�$d/q('��Fr���u6@�";�����\�F;�����Y���&G弒�������/�{35}9s�;޷�s����UNy�#�MJcFV]e�,�Q'a�Oj��I���2�X_�I���y�U\�͏+�>A<�0��q\c�LiK��+����P��0�≪n]�
,�Y�;�՘ J�� g���y���}��t=���9�f��q��(0�0�s��^�z���nFÖ��Dz����'��=g�E�I��s�~�4LEAj�p��V˂J<����.����YM,�{�HC�҂fg�Ko�Ue�OL��EgDrG'��S)��],��O�U��t��ɴ�$5TH߱.�[VT7�e��Ιb�� ���ZZO�s&-EZHy�?�m��Rߣ\�U3�N��I{�sEqЙ:)jh:Y�����+
UR�X ()u�Vqv���`��:�5�yv��2 �C�}��U��u�Y�A����^df<�F���UL�����@�
�9�	0	��)�k����·�0 x��s��a.��ro����?̮U!sȂ�p`�P9��&�~^�"��K����84��J�o�/!j��f���c��
���1�ӑּ� U�O�||�M�U�jv"ث@��Se�/?e�eK0d�K��P���-EA���c�m�X�=��A�p��/ah��T���L	�*��2~�2���N�a{��eLΤ�$jC2^h�>��h�l���;#GӼ� <J�إ:U���b1L�f8Zwfc�u�\ט�C�ܣ��k���.��7()����f�s��k�����m�e�V�x/��K��~MB#1W�.�2pZ���t\���%W&��vb�o��x$v�	��$V�螖�aSݲ;W|]P�~̭����j{w��ؑo߷��}e�B�L�wS����${�|F��@|`i	v7�+�ٽ��m�+��q������R���xi6E"��@��I>��b�i�hC
����E��g�dx��['0$��͉�b�R�}I�m���f����-3$O�:��l-��2F���@5��Ğ�@,�V9�C�(!�T���#a��M2�򊞚RJkq��B��ҋ M�$�3w5�g�/�J�A��5�g�PO�a#��x�
v��e_�951c�$x.
;)�Ac�Ƞv4;����+���y�]���D����n{u&�;�&��]�Pu��w�SdP�p�r��B�dd����h�֌a�~����8�����Q$V��ĹH�`~����ߛˠ]����h�N�4�fCK�����D=XtD=��Կ�-�qܬ6غ^�?��ڐ����x���3����h;
35.�g��E��H��HD��^|A.N<4'�H3P���� ���������[��?Jgq����%$ɑ������j*�!�گ�����v�'���L0���F�/��<�h>(���� H��E�jz$�|��>�RU_L�RuCNFo�a��(T�-��Ė8��կ���Wu�.FҸ�����s���_��>qh�������g����_mx�x�i�>��4�X�倶5t,��������^��u�.OhS�2���i�^�6'�����ܶwߏpܹ�˄���[�r�So��Y��0X6���=G�|v��*�R�����I�nL%^��7����Y�J-Y���t}p��>�����'hm' ~\eϊ�^`��h(��퇣�~� ��pe���R~�o[s��N��b���\Gײކ@J��▪�<OL��)΁�����d��^n�7�*\Qhi��AT ��G�E����ֿՁ�D�}-�YQ��w�<li2�������\��<>��������?&k��Ŀ��\+������p�����Ӌɪ�L�E騦Ƅ-ϗ�XE�9�)Vd��_:<9�n�jYyӎ8��D�aF��"�w����`q�_�76���Naqqw�Uf>�Q���:��>�:�Q���Z�Da���?��ݿRܚ�����,����4�m�4��&�y����Af�D��S;��=p��M.D�j柀�	�̶Fŧ.�xVf4.z�{m�5����*pЯbɄo[9�?Z�#�� cv����t��X�l�B_��$U[E�@i������˄���-����u�L� *tj0�t\�\��T�j2{F�_J����_o�+�ܨl,(-�ը'����j4r�h��;E���Q�`����:�g���I��5�̎��R�Nf�KR/Τ+��7���«V0�<5��?�L�)@�O�%1�L~�n���Da��5G|<!C΁�>���Al\o��eq�����8$|^�4}
���[Ȼ�Pݹ��!TQX����?͗�Z��qK�э- FV3��<����]��Ep��dR�zRƬ��`�����c�@�8�g}(
�6G&;z#�N��JҤ����C�GҖ�<P�����mvEM��h�vf�!$f|�4V�k`J�O�ak�������"���di���#�`���$L����V8�1�x�tq�e}� p�w^&/g���sgb���A�k�^CC���>�������/#oH� ԯ�.XCX9ձĜ�ҮcB�[;�u&:VWvQ=��T��6_Z)��Sx!�����k�6cf�Aѿ̤俾$�A�$P�ͩ% #���*v���N�����Xʆ�ׇs��M���${�q *��˵��.~��4#F��ev��u�'�F�a�AO�]���+�~���m�VU>�ԏ�|���#-VCQ<�usE�)��Q=�h�vM<��ZO�7|p��շ�xA`�?!�9�5A\;^C����X@�:(9�h�7�V�P��;���܇��0�������K�<OX�s}�����T^u��p��g0�,3�5���ڭ��h����b�,TC��i(/�����1f@"I�������S��a���є��~��08E{����pi=+�@��ngø�X����%��S���#A�[�&��<lŖ:�N��'�rlH|k�;���Q�c�����a!�`AfZ���8��޳��1��s����h�w� ��͝X���:.�����yi*��(�x��9F�����Z����E�,<��'�
���U�6A����K!�d�ʶ�Xخi;Q�dbن��%�ځ���2eui� $~��c{�p:h�\�(s�+V��Izێ9��j2a;S�����q�����^�=F�O�j��K�1����H%��[5x뺦������i�4�9��//u�[K��MӝÏ���p��SfS|I<;��6��c����j'�1`/+T�r��8�=)�E�L��ZT�s�s�k}�=����;u�-�����hB{����FY*�mR��LW@{��ܬ*dqI`s���,����n�:��el;�	��0jI������O�7O
�z����}ʡ	6���]L\����וX�"ه\�~�<h���L��6��Fb�&��&�d�7��)�9�p���q�b8C�;O��5�ƺ@r��^�[F#�]�ٱ�C� kcvyS�W�M/r}���)q�N��\�z�#��_�?�o`w��9(VN����L8���1������':)R/I�b����^xMS����#"~ֻ
W���!�:Rfԣ�0Z���įJG�TvW�']*n!Ig4
;K�[n�V�b`��ܝ���"��|��E�SU��;޲�Y�7ޝ]���+�Ol����Qr��݀R��8|���ݧ�[d��Xϵ���n����;������i-��OJ�T��]P�J�#����|�͂�4�[?)"�i��<�ز���S��[O�?:���P����&�O݇��IL��Ȫ�`!�v�,��>�%����Q��~`t\1*+�D�+�Z.�_7�!��f� �~��b�u3�G\|��dOB�w~��nX�"j�U����?`�BZ�ZlRD��"5g�9Jm�O��E�߷��bK��b�>g� ~r.���ɤ:5�e_x�ɻ�=<�$���s0���p��:7[-n�e�|�k��u}Þ��϶o�V
�7R���}�8T�)
�oQ�[�����Ր*�
Cdv�~���ᦌ�2J�_ً���x�ȬvA���I--:�9�7���׬�hw[��0`��M/J��c��y��ªOx<� �/����N{��4�A+���߬��ќs���3�y:��=m�1q�dш��&Cqb�W��̉}���-��	��9�R�I���;�f�}�b��Rr�>�+�2
\���i� ���7���i��Y�����tՉKn�����n��]@+�����w=H3�У�r ��ǰ �x�0����s�@�TcѲԙ*3Y?�߯�q(���J��U��ڞ+2����2@��o�|(���p	�L���<[-e�)AG\��j��m�
U�8�=��q&f�����;l����i fn���=q���z� Q�3�U�����p��t֑���"�1�Ѝ|���gaVu��WjKK�P������+h'9b��x��>�)�ᚭ�_�Q�A�F���P��]~sꟙ��"u�Ғ$�-��8� �D�˃�q[[�*|N<Ń��>���=��\��ن�+n�Q��$=Q�l��6c�fx-��5�c�/ZNbh�09湼�e$��ߎ��I��!�B}��4�cK�Ad�UzO�+Fc�=Zu�����ʝx/�UjZ-��i	*H�Y]0'܉�yY���L���SPi�>2h�o�v�QH��	�ԟ!�Wq���8��:À�X2&�pS����f.��0������1,�& S�a�XE�Cμ��ڍ�ƶ�b���R&Z��A+�e^c�Iy\���p	�z<$�[���zH�����`G�B,/�UP��V�]�������k��Թ�!e�&��{�1�%i,�9(P�V��Z?W��h��N�<]������5곔?���
������'\̷=;7��'Nc��4R�E�*�!��~:��B�
�:����d��'�l������k��l
>���T'�׃�%���c�m3=X��� u����372�q��-0D�[� �-]?�oz�;�:�ƖG\^kCJ�l��.XA#���Ǐ�`��9˝{�o�>��'3C�����T�0�0�\��:����&GAG��n��_�]9j|��@�l=PUw�(w�%�J7�)"�ξ�Qk>
+��I,�����#���8��Oڶ �C\�qᖒ6��M���VN�g�U�B����,j`�!��Ĳ˃Dg�Z�?���~��(���dm����5�y=�[2��CK��'��N!��g(�1]٥2�,^f%��)n)[��z{�n!�!��X�Uy�5C��� ���b�V٢5�2�wu�u�����
j�����R��t���U#t;X�b_4vD&7�"s"�1�m����h��e�j.���a}Fpl�h�bEh4Cb7bNl��.������Fwт�d��ږ�,���P��s�-)�������z ���v�����9�����Xb%�@�+�;�D�3�B�+�]���<E������� zק���ސ�bM�ʏmM��2�'O�K�L�����q���`�:�Y|��_�cvU�ߡ�0f�c��ƶ�p�9�8��{�3t�л���-�ܞ�T��)�$L\;m�ҥ���O�u���Z��k����H�����	�
S�ѹA�_΢~����/}�,�5�$�$�}�Ç]┙m	�س�|�K�-�{����~0"#�o�;�ucųxD:B>,��a�[�W�7��O�1l4��b\�V���)��$�9e�'�� <r�y�PV�
wAI����/�+���P3�ED���5��Ա��ͻe�:`D�d�/o~�,�$F�3:�J�6U��e�0���kþ���Xk�6�og4�@֚zOy��{"�Z�^��� �Oo��Ԗ�zn��g�	˅�<��S�[� w�V��SHdfޛ�U�B�j��C��.��O��7��t�Jc	�X	�°͍�#��/�D��vW��5��S�P���(.��]��U�G�w	���Fi��;��g{&��b4��b����޹H!ٳ�>a>�˚ʮ�~s�^E��	B"w�=6�W�v�ҭ��Y���8������9-��z���b�����/P8���Q��D��i�So۹ͣ~p�4���ds����g*5�N���2a�+BZ��5&s�6e���Έ�� Ԓ&�sx�M_�!�ur�]�9+���{����Q��3D�E��&'�g�dP��`�`��1����VF��{�T����b~eBz�JF�!���VbY�~AÂӏ�x�<�����n�����ʕ�r���k�h�G��ȣ�ؓi�����
V��,�ɺ#�b�5V�=��#7�F���3K�t3�#
k66����Y�s9�m���J�^��f��qQ��_?B�*�e��2ʸ����V&d�����ا�qU���������Ery��&��r?J"xT�~"Ż�?�FSd��JÂ����}�S�F���SF���PI3*s.�������Č�z(�]Y��Hd&`� �jM1J�;�pJ��/ ���ge���+3�c�̙S�d�-?��A��%q�� 8�۾�n��DԶ�)�1g+Z��6���_FL+�e0��b�ᵧ��Z�1T�x`��Q��7����ӬH���e6!��l���5�(jޝ��\���9������Ўg�)�py�E�I�jS�#م��htҙ���@�&]OUPO���ul�Rn@.Y��� ��)��EA2����	�s�2o�ie�*�|	�7@ip{�I{
���k���(/���� 8�$׼�C�&�������P����w�_#�S��VS��q�<`N�Z�N�Wl���I��qN��C�#(X�/������s���EU�����F�kU��o;P��E  �Oܬ��TLAܖ�ȍ���g��O�LSi����u���!��)n��RM��8�sM�d��y*��>�!]D�s�H��P��I:Qv&������Qӗo�e`��E�2��5u�#=�J��pc�eX�������Zɡ��{Gu��f�;�3�ML��W%|^3�rٕ�N����j.2/k�A=TT��m��$�4�f��7Mh�w���_Q���C4^Z�'�gʏ���,Qt�������sQ�I>(�B���tJ#�O<(raJ���~��S�5�Y<o�������������>X��?�4��R5�_$�4T���e3�]�:tp��D=���~��m=�,^�������@�A\nMe�q�W���Jq���)r�\򣺮���8к�T�d1C�r��V|.��)QA�6z��jvM��Kk)�����G��f9V�i�� �2]�i�����l���aĹ},�A\��ä��
8:#���=cb��\�|HÂ�:�c���8��`΅p7����:�K��e-zJ�|�AcI��v8����[C����m�As{��4�ۡ�~]`����ȽM@>�/����`&k��P�W��l�@�,?�͇��h).�?Ag?���Z��츈�>G�𻿑0,�Z)�K�3���uីζYɰnɖ7��l��9j"�3M�?�f���$���]�q���^⍖�/�'԰���&��s�� �i���_��=�i��9Ǧ��n�#u�N���-�з�V�'�ķZEs�����*�꜒���zd���"��K7�!h���ܔ*����1:�i��_6�MT�i�>J���3eȶg.�w�%-��)p#J��y�?��A�7yU΅BG Q��f��=����6�C�Y���Ϣ�^��J���]��錰�pFk��DU�ع9XİR�T��H㽌=#����$���q�*������d����œ{;�����+Mഋ�P%�}�u�3W�"D����L�Ɩ��x�0Q�PG�b��2v�?|ܬkq����v+�D��Ygx�gH�Ȋ[z�&�O��I?\���j�K�5��9&j��B�;}�a�f�Q�Ms#�'0�HJ�߶�m�9�N9?k�x4�:���X���
�11W~��6�JhD����|X{aَ���^8�ṕ��z*���K'^2c�[�X��'�.'l�v�� ؐ�)�g/K���A������t�[������̄��"(G{�e�b@�}�=tk3��`ʂ��}�LEx8_������ރ3K�#��V	u�]̄�܆Q�y��]���(�GS�	XI���'��$a?����U�S��g���u�����MZ?i_�z�p��G�2Y��$�b}>�U*u9r�_�m�z��(K��1�n
,�^M�՟0}�������xw�KCLI����;TL���Kt^�d�u�YT����I(Z77��x�CJ�8gg�Ը?������/�X��a�2�D��
N��SF���'d�(`T�3��u����K��)q�8Q �U�W�5*@x�n����6;��C�N#XC�#��������2t�H�ֹ(V�+��vʃeU����č�r8E�I�l�{S��� ��H����ڭh�OB{B��r�캗8����Eq��)��tc䖺���n�!Qe��G�:���̬��#�d�-D�3c*����*b>��X�p`�׎�~?�B���Ei'q5�h�,gJƚ�տ	�0��-��W�)�xn�!������o�^��#�cq9���ɪ�`h�H3��.}o O٣o�0��k�(���eN�~ߙﾆ����F�Z�}�6`��O��#�sW�O��R?�R���Y�t�t;q�-��N1���N �||���c���������[����#}�8)Nu1.��4��qs�
�a���:���}�9����x��۵��,�D?er-���<@�Mc�x��6��Lxq���#��0��0$�֕\�(�c�"��t�P�G?�w�Q�E\�=���QC#��w*�� ���eq� ��IH����/ /,��.�� �K�v&�u�C7vW�Mʮ֚����;������7JE���>x��}yGh�c��l��j��l&�/|����$�^{�1�0�kc^���m��}߸�c�e���c �d��y�L� ��%|`�@�t�Q����ޔ��!��I�3�y���y[*�	�$`�h��7Y�J]E��BP1⎷��BC*dFV�E�@I��~���]?���aa�Kk�4�J�s���,(��)8ބp�;,-�W��Kx���		�%G����F��Xxu_HJ�������<Hy㡻�;�y��o+D�R2�fB����w t�f+E/ng��m0F�z�1�fЄ[gv�~�%�X�
�˓}w/�g�y"�\��r���9�B����&F�����U�0\��.Ͽ�0@#�ߒ�Xwk&R��:A	�pf;�ba����p�D�>�B���3�*�$��2��
�Vo4����q�8���Դ��5��1����W�K�أ�F�ѫ��2�*}�� ސ��ؗ5]K�l��WĜ���ŕ���1l���ЙRK��j��3�l̕fϑ�@��8��6����Ȩ8Z:Ŧ�|G�s�����l�<i�t��.���?�~!�V�8-�uz��t7��ֈ?�U�FZ]b	�O �1^����&�9Ac��.z�jUjZ?I�C��J����X�8%�n�#x �B<�a\wVWmԒ:"ev%Y6��,��E=Gd���Y. ����A�<*Wa癊�х����a=�K\{��b�J9&�ݾ�I�c��kG�"2���0D1V$I�G*�e�Z9������\�O� �p�,�Ѿ�[�:�t��Ċ�;��e�g�G�XGfoh��?$nDE�E^­��i�j��u�����i�.��t�דSw�y�;#��+W�7	�s��	G����F2��W@V���
��NVu�oIe'���"`���6(k'tI������$��tnT���J�'�&J����Co+�QX���w�`F֜fq�]kU��;�G!c7����yb���� ��N[1̥�V�B)ڑ$�@3w�AqR��~��dK��'�Բ�7�q�ƚ�,�����]��w�z����# �0���l�W��΀����ch=�r�;?߲���>�e���"�m+��Ǡ�w]jF�lU�e�
]�Y8� �,W�	�	�y�p�2Y2.��E���<�,�p[��+��Xƅ7Ԛ������"x���I�|Ed35>��<;0d^���K^�	��d��3U?��Nf���o��x�i�K o�~�=.+K��u������G�p���)3�;���3��N/�	H��H�h�������O�KV:.�Yf�z7���y�<:��av'{���ճ�E�X�Gdg�zOq�kc��+��=���5�X�{�B"�
��R��'�X�__Ϝ�}�u����ƨ)�E��Cq��@<c�5>#l�>��D���'{��� �xe��b/� �D�|!���,6����E�rs����KꐂmP� U���~��_�t))G?�&��,���ߝb+���YJ�c�B��LSIyX|<i�(��G�����t *��px�
+]�my^�~Mo��B{����ƈߚ�n����Mk��y����&����f\��"U#�.�"�`T�
o��FJ���^�Zw�V���5���\�!'0��٠j3a��1�����F�[�n�i�E���G�*ݵy�O����0y��CW��h|�e���3;' ��]ڎ�"k��{�%p|����E�~��l��#\�<�B�������:c�>�mv������
���+�V_l�Wa�*�]Z�S���v95	F�V�Bܓ_3)9}9A�z���+m��ν��'Y���H�� Nܦ����]���K�~�&uZ<^�"�sW8Z���Uz���uf���b{�]�V��D�OZ�_i:��5�a��:�u���l[��	�&���/�>�Q
��K�e���2;i�^�{� P�N^�+�2J��4���.;0)��K�cSMz��!�d����4gZ��+ç��J-(�{��Bь���^zU��Ű��}j�5���R�?�Fnq�=o~�]��oQ)�:`VT{P�M����I49��
UN�o�Z(�/�k��@v��p@^�>��,���*�eX�e`4�3
�w.j�x(xͨ�����)+�˔�����Ua��|l	_$�hU�X�n_[J�E��b�F�%�L�sv�X�o�t#�7AhLid�<��H�^�+�������6�H��%��V���:͞����p�@�3}�i�8ǫpq�)�A��p�p���v�o(���6qx�߲$�HN����R��f�>^��O)ɡ%�)3�}��������XO��J��E������5pt�mE�E�����aԊ�\���7��	u0��}6��42�T0^'�%U��*c6IM���r.L����D̐�֍�N_�f���f����G"aw��pRO)�Z�L%��t��v�7'^��qgj���F�����x`&��n�ň��6Wo����v�o�6?w�z)�Շz�\H#�A­4[-� ht�ء�e%-r�k��B��I��*�|��0��������.:��WG�R���l��3��6V�kR-6��~@GYe,\�ht�M,rT�jE+����рˠ����wK��8���C�P�G�Ռb�:�
'��;��<��W�ЮHyXw�[^~>�p�1.��L>�p����b�%�]�����T9�L�K�'��.���?i1^��^*ۛ3֔��#}c�Y��_�����j�.��t����m�{���O�R(�g���3�4`L��,�~+~�Y�~�n/�+�c�+h����N�+z�7��n�&3�;<@�L�xl���/$K:d��q,�:R�R��������� K�LQ��ꎳ�NQ��p�0o4) ����(���)���b��us�2m���*t�Q)K��E�)�:�S�6)��f�l���R)��ʾR� ���|ՌU��8@ڹ�0��4�)Zb��4U�F�����ݝ���&]]G�#:\�5UX�yG�3�(|�+��E��of�_�F��.��7@m,����$3'_�P���ӓַ�d]ܢ<g.�?!۷����K�tAe����������F�)+���p�����๳���5�ZwH�o�Y�;#F,�*kz֨�,���P���͈є�
�V�A�f|g��WM���pQD��ߍIrm2,Ɗ֫9,dgu���;�hMq��-� �v�]��0�r�>`�|7���U�_6B^6�	C��~�Nڔ���D�>f�k�龒�Hw�/*e�\���=Z��%��Nq��8���c����`�"����r���>zv6��3#��D���eʖu�ODU�TN��dP��k>&�[f�a��>N#*eH��NbX>��F
(.��5Y�{�ȼ�Sܕ[F��
ٟZ:�#ڻ��!��J�3��J�S����*|O� �X񰳄�"6�^C���I��	м���9���?��������eg-��d������6�=P��rr\�@˵�����=\Q���;҉u��5/�W����K;�+�f\U<Z`�OR~F?�a�#�n�Pj��R!Ds~ �Q:�v�ރ����%�?~1���ae��*b�`z @HG��@��}��d����������b}:���e{g]��UW�����Nd NW�;LZ�_�o1L��	���\iͻ7q;z������@!ZϹ�	�!��HB�LQ;Ba -����[5f�~��W�F���_��^Pk����Xx5.��ʸ�!8����HƍL5�bZg����H7^,�!ə��P��g{��I]o�	TD����yRϦ��^U��Pן���u�P�Z.!��F)s���W�)��u���g�.eEt!�ʘcD�Ik6pԪ��?�;G�q5������������I���ֺ�׻�W����D�������W���R�F�:�U�Y�n�z��X���R�eDx����dYJ�)@��1ϡ�_CY�߾�:����b鉜�ibf�@L�
'�t��II�ǯ��}���Dp0a��0��M�ܔ6�hת��et�3�%!�m_����?Aв`����ɕ������7�	�ɾ�O��b�Ay<��A�D���"5�[W���{}��&��t_�f�nш#��T���h��`]����g:'WL�~��M8��2���n������e��nԎ/�sM{Q �bHL)���,�iS7Z޾"�?Mk��){�TД���#r7D5\g
�,7ٷ�3dUi�-#~LR��R|��cV�����Ud ��8�)bz ���SUz��B/nw���'���F4w�ut�������I���ˇ���S�WŌ4���c�âx(�\MZ�ӻ���L纣4�.���O�g�,��'���]bɛ�>H7����m�'��3���Rg��߉�2/��J�S�?�K%[�
>�NN��Z��!+��Ǚ���3.ll��:C�>P��SO��h�=	����@�c�Q�MЃDP$���ՙEb�OHa Z8�!���}/ ����ђ}���d� ��r����M")�.��ru�ß�V��|��^�1&�t]$X1��k���X.���<S���-ڲ�BD�Q����2)q�^?0�-�2S`K�ux����s�7�aJb8����&���W��������b�޾hS�#c�@����+Cʃ�t����Bmۜ ��w��b ՈN<˒pg�4Hi_�- �]��u���WQ�O�~LQ�&$dӊ��b�~���`�O1�Xא�^{�<@�Q3Ϳ�>c�x�~�Q���(d�N$����xG$�Ӑg{�w9� �5s[�6���65w����par5�������}�[Y���+����_ח��*G[���vWd�ʷ�z�dԗ��t�Z��d�i
�C̛�2cX����c��ڑ� ��-�-�\�S+�o�7�!�c Yd�s�Z5��Xe�&M0�U���G���	�}����d�'��#KX�|94t|�Z���{uF�g=�
��F�6��d�����ZDb<o}�Pr��MQK��-�Ч?_���o�3n����J�Uh��.����뙓�L4�<d�;NL��%��e�6M1 �9�u���"T _�[�(�%��9�6�&�x����jBv��G�L�2:g������ߙ��)O	#�q1���[�
�`C���`A ��W���\��z�z�|h��Qs��v�w7s�������sG��CI��v�4@�]�\�U[�$+_�(*��q�����ܱ��g�h[������Mg��Ə[�~�ɔB��z#b�����&��n�Ԋ�F����j̛�ʣf����j�E�.[�>���#��1U�s6�c���鄅�w�7`B��¡PQ��<o@&���o<G����\G�eRm7���5��v?�X�qg�����g	줕آߌ�f������d,�� ��n��t=d��s�m�%� ݸ@�d�`�
Q����
,����T��ԛ5Ɓ��m���omy_�$[M��y�S���yJ�{���c_�6B��.�7��⥹�\�v>K�;j���	PM �v��p-?��<� $�����U@�e]p�M�m,I�HCaҤ-��ϋ���@e?:7��}5X�L���3x �2�_��(�ceAw�j���a��b�^��p��C��&�
r
l�[ �XL�dXV�_S�[N�ւ�z�^0"�N���
�H�H�0Q���p����~��i������E� ����y����3���J6��nw?�&af��f!��v=i�\ESZv��+����LЋ�mv�u���t�@U�.���� �:�,��ы�d�����.��U{��3����)�)�ڶ �r�G�70�c!�v�͒S�͝`���@�J��^�쓓'>�)�-���1��Ɓ�OS�	��$�@�/�:�֗��#X�����*��DQt��M�k*;�8��B��$��T�o!��%������5�I�@���z��dBW���,��o�וAX���/��wGW�QX����Po XHСꤾ�'�p\wE�D%ld]����SJ�HE��v%��A�d	��op��A&9m\��<,�C�ZRra�C#�ylsV��~Qy�vx��Ҥˊt��V�,�&��ZJ2�O��߼�3�����0�"R�� u���MY�J�t��ϾDP�Lm"cr���ϔjK�p/L�����߽��ك����}�	�}�s7I�i3zu#	@F2}��G�EL[R�^��9f�(�5-7�|U�g��ғ-]?ӳ�<��Ǎ�/�Q�4S�:��	?AR"p�ز��1�U))�g����^cƪ��E��6�e���UBPS�LF��êed��wK�􃣕���36c�\}��۲��(�,�eٷ=�S-�#M�"ˮ齥��f������v@�������c��Ɠ�t�b}���ވ>aB�����cG�0���&�
�٬��3�sdCk��_��BI��$R? �ğ!���Е�c�k�����h����H�h�:�e���?cg�弻hƘ�����B�*��N?�еđ���ŒT�=b����Uq��A�&�b8+�(cr�:�����S(�x��Z~רK�Ei9Wr!H��9�W$�3(�:�Y�]��� �92*���r�ݩ	3ǎ;F�Λ�N��n����7��(_;f�w�+w%^h�S��*a&a��~
&�O�Q�N?�KK�*�C��D�
�jI57 CɌ�ё�#8�ؚE�έN��� 9��x����<�0�g|&"ͧP�;�x�?�nM�e�$?Zs$|�@����L��N>i���庡��9mH�6�8iXqIƧ���1��dO*����8����{���9ST���VA̡)�3˷��*�+U�A����;�?e�e���,�1���x�Di�X�r�ng���AK�I�:��K�j�3���#����xW�Nzr�,�%w��H����4 �Q Q�*��¢��^s�:�Ǧ*� �����52b	���Q�}�-"�U�����H��gc�n�nk��L�Ela3/�Z��گ�OA���G��x��Q)[�Ei�����|�Y;��n�G\��C�g��E�u��g�y���/��(�Q�P�9���o�S����^K� )`���la����1��Ov�@�к�L	ݨ7>�r)�m{_��Y�lBA��Ķ���S�hI�q
w#xm��3�5��M�ҝ�1�_2D�J�>����J4�I<ˀE]"���=�����[&�
���*�A�پP���ES��9N�;�绗� 9N��sK���6_\��KIY�
���!�s�g�+�F���f�$1Tl�>_�Q���LFq��"�(�J���;�(K!%l�
)N\'jjGX��Хs��CV��ie�nw(��fǺH	����q����q �R==!��;�q�昷�ﳪ�Buy�y�:���֟C�+lY���d����t$:���t���K���t��v�4�`�+M=A �}��/$�;4��zDf�+�s�������i�mtU�#tY_�տ�9-��UʠHjRo�������hM��"�_=�` �d+X��Nˀ1�5u\�i�H[�t��(s�Y?UHy9���n����s[�4�$��?�1Q��77���q��IT����Q��cG�ά�G���e)������t�mH�3�������;��#�m`�٘����=K�-�Q�D~�Ġ����޲�\E-���d�i�k-��l���*�-4����,v~��U��3�~ɀ��>�>�؏���d���2�Zn��y: ��|�c���,�0A­�t��y��Q�L�;vo=GR�A�/}>��`]�L����mk�}G�ߌ��we]咠��U]S�ݺ[�Z�����v���/} ��~ ��]S�2+�}�8��;�Zy���Ar�͵�'x�٫�WU�h������%@����iԾaB�8K�p��P5q럂�I�B�SL:�=~�V-.4�^����1Y��#)&V3��)m��e�Lv�E�fV� k60<��}��)�2[(�+a����jv��Ǖuo��+*�^#<�RR��!�M��~l�
� ��a�#ȀZ>t��QG]Tun�nڞ���[�lP<�����gk�>�3���9�1C�7_��`����`������U� �3�	�q͎������t�w�ӑ|�/�߅���f�N������A��@��4^���u��K���d��׽;8�?��N��;�I\���Δ��2bӁ����3��ޚ���
�ϰ�M�K!P�-�wL�a�s3;B�c8��<��7�|؈HQ�q�7�����r�1�OJ3dI/��^΃~痞@W��޴̔3qm�4R�.fgxM�
�lڛ,�o��@Ј�woĸ�i�f}��jl�`iT�̄��ʭ��^�+޵��K�w��z�xJ�}�d���������N�BGͱ�Ч:�2����w��nC���X��[܉I
����R���30������dx�$`(�/�R\'�r��@�ș�`����kn�Qj0��[u^S�l-����FBn�G�4��a������B��-r�ĳ.����{m�^�P�0�h|^��R�ۡ�AA���e`��,��$�V^�嵚
w��ko��ON��(��5]8��uE�&*�87�ӹ@���]���.�A;���^#�!t�5��}��{�_ym����P�9w{�;�`����:�������ԭ_?�E�L٩�k߰2��k�!����+jHV(��f���6�P�0�Iy��kR�OR����-Q����W��P����}Ֆ��H�E��$\4�Z�5U�zQ�x�����Vv\���Z)U��*BV�ТXZ�L���#L��1���ɭ$��W`]�5�2$)ݱ��A�O�U��k?0�%AǑj1�k y�u�ش'bZ��_iNS�L����Oő&�Leԇ��n������E�Cދ_z˳�@�3��8,�s+~/�?���/��0-FT��%@���Uj�~�Ub��2g��5����Q�V�;�?����͸��B�W�R'h�ܠϘɻU�(�Hk�B;��k;�y�]/ο�ۙڝsXS�R�w$�J�O`�b�aO�lm�Ϩk�d��8h�Wx�Vć��I��,nٴ���@Ȇ�ح��JʹQ�?�.�Ӆ�Փ�'���Z]B��^���vcp�)
��Q�������A�S��L��H��lyf'+���}v����
q�Uj��6$e�)�82���a��k#��C��,�g?�#�JQ]7����&u�n����P���?���ccr�&J��p�J����������z� %�7�|7@�����P��0��1�&�_��Ӟ.U�M䣯����j�^!Y� ��߼m~������͞����T�{*����Cn�?,6�7����������+xT�3W#�U]Nl���������ZŇ>1�cO��(:�$�@���r[($Yˈ{�C�(���ZĀb�'��� �b�]�AΓ|���>���]ۇ$`}��oj��.j�F���xa��Y`�Y��f��VŃ_o�]�/iv7�������'�$l�	�(���9�C�A�dc���.\�.Vzk�h�q����t����d�6����{�d	�Cm�kpq��bO��9)��[�N�� FJ�hJڤu����4�ɇ���,Qث��f^��÷�-���`�k?0�t_�X��(-�&6�+r�"a��b�u�����ޱ���/� {s���H��h�X1�#���E�AP��E\-�9�K�;��X�A�/��Y.P�7�vMϺ�|𞻚4.����\�ps<���QT�ı-�W�e�i")h�A�����%O�'��R��c����5U��@Rw4"�h��	�������8
6T���b��,pb^�B�Q��׳�#�5�ݨB,oΐ��&r�3�R��<U-h$����� `CX�i��pxn�0�?Nb�a��A/ª5�;[xsY*��W��X�.S��%��Cq�u8��#Z���w?��j�HEV�ir�E�X2��9����o�r*G�w�>Q4�x��k5e�l1��3�;��4qn����/Ceȍn�m1I�Np�t>��	��8P�G8n=:��
��>Ұ��Ē���o8���7�^D#f՛���<�'��(�NM|���Ȃ��E������2��K0Zq�l�m,R߃{ʯD�=���$�k� �
u��O_����.�~���ی
5��X�����%H��>�����`WD_��4܊��L|��@^1�h6:?
�'O1��P�Ϭ6���앛�����j ��%�%��Zs�Z\��_p��Y��0#�b�����#�
���
�TmW'f�Hy���*8��,��	[x��b(�U�3;��.�K��֋�rbo�ݟ�-C5�?��ˁd����Ҡƍ;^^��0:��{%��	���m#M�:��ao���e�C��!�/�����V�X,P�b���,��
W�"S:��l�@�����7�P�G ~��H��k�mtvK�:���#�v��,$].�g�^�#Lt����8U�F��-�ƀ��gX����+j���{�<��0�4��9�JB	�P��A��*��0K��E�\�����;Gi���+T_�L�I���A�>�� =�
,��C���O�a�M����N#^���� ��$�cԀ!�����y�s�N�I/.X�X���x�\����'���U2�k���%�段�Q�� ���*�G(pU��g.x�	��՝���t�� 	;r;	�����o�P���߿��8���m�b��yK�I�+�~����n��D����^�e)����I���N~�
�8|l�F `�È5����� ���0�#���P���Y�Eܫ7r�� m1a���=4��C�˙�	JXF!}y2�S��]�7w�. 6�p+9J��Z��j�Jz��aX�Ǉ߲fk�5����Pոȟ����Ӟ����Qًe\���
��~�����Ⱦ�Vh�J�媡��%��|��˚�-Di�E�lo{�Љ�o��tP�q���;�y"�-_�YF�#~�F(u-���h�$RQ�9Lfz�B�L�9[G��m�4FO��*�u��tz4��n�ǫ}�*��;�c�݊4���MP�-/`�ԥ�}g��$K`P*�6��x��z�9��H�>ݎ�ٹ܊1lm���s��I�JV�S�i�=�`Feڝ�5��wL�E�w��[��J�xT�LP�"�`���M����A��J,Q�ϥ:���8I�{������_�7VH�5���-��W{�� ����:}�t�t�[�`�j��-P�N���	�E�"cTaP#ɆDT�s (̋�
G�N�!�ɐ�t�X�Kt,|"^,�9Ly,:qA��9r5ƃ�$-A�@�J����6��}sRs� M�+;��;�.�"��? ��S�'��q�K�>g��P�� ����b��T�
:��|L^	V�#�wˀ�S�=j}�,��eՂH���,�k@"G}N������M��Eo��N��c��z8�����vL w��1S�P�^tn�윇����Qv�f{�!şI3���}�����J$�)[v�ilhu�����ÿ�b�;�����c{�����j�/��O#�T<���D��	�f�,��8~�زq�['����ŚA���MM.�k%�Gj8EVܚ	����eE5Xʇ!�b��������2A���fӵ��v����A�5L_,lKi��hr��T�v��?k�^� �g"jvE]ʔ�%�z�ekZ�fӟ\�Ծ�*��C���n�R��(`����چ��|���C�$T�ΧS��i�څ��e����l+S�y�-�{����XK�B���ޞ.�<>���:�M*��M�n����L�MC0Hso��X7�7�`�duQA�$Y
���@�O-U�x!�\*Slz�5�{Ȑ-4G��̂y�RrNL�N=yd"PǱ$�y,k]���K����}�,Q� ��R�q���{��Ή&^y×~'�]���<,�H�~�
P�G5�œ� JY3rl��6�q!Q�~�&�s���[��ث�&a�MY��a�S��&ۥ*�B��D����B��vۂTgY�y���)��
�
 w�_�s\�3�S�ۨ��N���� ���	;2��)��?�S����.n5�R�?�O=�2��8���+�S;|Xq�^��/�kp���7���x��75�D�;��^N���v�~��d�^W�x��� ���q���b#�e�k���VZ��.���~WK�|?����p5�>(�V��I����/�F��V̠a�s7�І��\ڡ'[�%Ŗ�^5�%~��`yA���UT�ļ�[SG����?���W�<�K"X�- �D2U*�L窔�n���*�<�<ɑ�lb|�1�cl���!Mި3��V3\�����>%��
e�������E���l�?8x;�O�]��4r�]�ǻ��iM����_�1���٪X"�}����W��J��gS]�`ϳ��b\��6���8� ��u�7�r�%I<&T�{-ta����=å����aO�|$Y�Τ���8[�q�4˼���st�傧 �T.�J�(��i9\�����B�¼CBJ��Sj}�,�n�陳(�ڠ����B%9Y���74��KU����{P���K�2��C;��R7^��ZJ�g�IptC^Z ���2�u2?�{~�W����-	iS�?�f�*����<��|�>֎�d��7#�[����7Jng4����Y��}��=㈐t�����s_��f��~��_Mt������'�(\��B{ܚ��ޤ���X�[��]�L�����8.����D�/L�@������k�*���M���-��A&�֒��F��|�q�3$�W�5f'�QP�@�<$�mk�CG�r�H�33���JC)�4��i��J|D ��%��:ü��$���j��P�-?��2���i�3��{�x��؁uHG B���e.~�r,kR7�e	p�ױk�F��P4�����K.KS�H�W�<"_u+��$F�4�npA�/Ϛ>6��\���˒H��^�����|�Л�9�2��Ceq�Rb� �g��3a�t�a�u��U�vMǕwW��xL��>%q�n�^���#h�@�򆼽n��O��$�<��c�X6�5m�z�S�0�:6O��)$d�
?��W6�Z�:S�4�^����v��a_h	̛��&b��L��V/;Xm�Κp.;.�x˳,}�e"�E��O��<�-m��t�zH�PNb�"8P`�*����9��̊�4(qi--n��m �=�6Y�����5��λcs�e��[g.;R�4e�3�r{��e�]�_0�Q�C�M�2zG�a��|�P�IX����5&B��#l-|��y��k���#yY��h�ė/�nc��x;�%��ϳ�1�K@[�����>|��1��aC[)�.&�|����:���s`���&�܁�V��BB�4[��{Z�bL�.N���YUF��0 �R�_�Fj�͉��˫�7��~57*�Ao�3E.)���b�f���R;��̺�}�A�x�t�7��Q���{r�U�s��ï"����)�6������6W��~�?\Pq���<َ!k��2Mg�G0�d<�/�~�u7J6�xk��V�jv�5q��D�\?��(!��j�1zw��b �8 H��m u�@��H���%��$���8�@�S@�I��->c�mV���1u�m䨯��];���Pj����Q�Rt�MJj�D��$�ܢ6�����ó:9RHjЩ���lr_<�5f|f� ���'հ�ǫ}xW���ȼԤ]mx�DH���`^��a8C���	��2J��ͩ5��-
����F������A ����6����3�����s�זB2�ӹ9��������ͥo،�9�ܑ�m�B�?4�7�g���c\Y���}=QT��C���$��]�6n���.
kg��t-R�Ѳ7��z����@d����(��B6�&�8v����'ք��]<���=�n��Ę�xlI)z`�Z�Q�y%^F���+@Y��(�js��ux���?i,��>���l�s.����X@�C�-�8�g��Ԁd����!r���r�B�0,g?�+0�]�([W��r���`���ȗ�W�W��!J���a�ivOQ�U-�K�RC���O}������.ڣ2�C� m�P�O���J�	@�ϒf���R��\���-���0�c���t��&|@: ��8M!/��[6M�ʯ>�ݟ���%Wx���!#k�Xj��m�i&��0rݼO_��2�1�����n��,9b�mÓI�%зf@;\M?V��I�Js����-S��:��1�lR�zy(�� �g�wG� g�f~�Hz���D��)02I%��0�(%ez�	e����(�2�&�}��g�1[r�TU���o��$I

@o�٩��7�[�PRȶW� �X.�m���zv�%[��E�)3t��i�t�O��
��x���<��p��h���5ȅ.W�?[9iN�_r�����}��N~�i�������z�v'��d�Q]n>��8u[k�9؎�e\���ءf��{�k���NR��V����%�OlA·�Vǡn7vu���� B�ILj-���nNw�,��ڎ I�5��p��N�� ��Z-(��-f)�]W�hK�Q�'W�w�&�+&U��[{zpg�OTz�5�؏u4�	�}G���41��T1x��!Ίr�Gw��֙�1�sx�ey��8�b�|Fk��.\C�ӎܻt�';�#�읤4��-��E����i�)dqG�M�Hb�������і��<9:��%F�كp���l�[^*����G��G�?N6\�Ҟ9��!ݭ=�t�l��,-�w��/�ܞV~z _�'��9=P���ϓ��1I%8�|9](�o���N�n�d��qT݂�Qrͤ ʐ'����"{�6�0��(Уԥ	�Zl�=\�W�!t���5Li�����\5�'�6چ-^�2e�D=�-qG�D��	
'B�Dd���|�&��t�l��/	i�u䱞�x�w&�@_���%�S��OI�n������{�U~nkD1�����YW-�C�0~ʫC���x>?���f)Sƹ@���pl�Y"��a �Ld���hPU�|�<���7E�����7���k�����X�����=��W�P�r����ͨ�շt��7xY�A�3�����us�=�3�1�������so@Y��~�98�}o��Qt�+�����ga��|j�K�IF�����ҁՎ�{�Y�2��Q��`ܥ-XGV�0gM�C3
G�}��]�I�����&�_�E6N�.x����M�o��N�#��5��k�Y��pq\f�	�J[Fx^<�E?L^5&�x1��/�����C@o`�x;�F��V������o��4�'un�����{�m��0�E�-C���\�ȏ϶ߩ�����~���(GJ,PZQ�+������Ξ񨒺�<��P����2\cu�zG�c+x���a��&��NP}�����p�,��M�������n������BH�u���(
��Z@�bQctc���	�B���W,��zܿ���ђ�wf*��.�!c5.�����f���������Z_Œ2�4D�m"���^i�m��=��7jS��V.2!�܎�f�LnM�ö���ݕ�\�d0�c�GqU+�ա5�>B8s�q:�LvA��
C����؇9���R ��>������<��G?j�~〚���Q���"��~�Ѡ�1@�"I�[�`�v�Ҙi�D�-1#���b@`;��G��&���o��������N��Z���[퍶�q��jΉi�m����ŗ`�Ru�5W�tJ����9IvIm�#'�V.��7�oX�����ؙ� ��0x�?�s�2��������N,���^ +�Ŵ�gjl��f��*�)�R6���h���[��N��_��Q��v�f���b�ԯns�8WB^�Rܡ�ϴ{��iJ���{q���G��K}B��dBCev<�[�us �&}�D�R�^עz8-(���Kw������6p��z�N��8y��K��8�,5w���k�q����UF�+m�e>�roN�e�i�* D�nc~-E�o�����l֧q�em��T���:IN�sϟ�M�Ọ#��{��{���Nà�I��7��N{�޵���6��y�A�/�����%��$�Z/�B�ȁ����@��Yc)zwrW������Þ��D��� �J!�c���b�i�I��t\�2<����<Q㈦��T�� be��
G"G���F�P�'粴����$�;�����}� �9%��h��f3�Y�԰6}���)0&q��!Jq+�:����?��Ǒ�PaN�@�s�f"[��2ώ)�%��T^i�n�|��숿�i-�pג�2S�6��OT_�����%.8�l���k�L(�ڳ0��|(�k§� Z�\��ǡS3�����T����c����K�X��:���2�������:͉���+H�|*�����C�d�S{f��� �d����&ӟø�&��Kӗr���ݘ��������ڤ���0z̭<@�b�����nK�n��0aG��`ۆ�taѺ�A2��t����0P_�����t��Э.��\ֲ�i��g]Ɂ��v��;�S�&į�#����%������/iʌM�s�Ǻ��vRx��,���	ru�w,��0�S��)!C���H�9�<�T����U�*P��ќT�
фǄƅi����?�(`�n�;�UCG�[�Pe��-��i3��p���6��wt�7YD� Dm��G*·*HEQ$0����53D�Px������q�����M���ĿJAu;F�ʓ���X��D*���HX���DݒsFw|���a��;�<�۫4��]^� ҂NYG�y�'f��<G~ͥ��9CՓ�����X����^�3!6,ULR=��[ܐ\�@L��/}��*;�'����v�J����:�IT���W�q�M�R�G�Qjz�W;�KfWs!�{\�����A�"WE�>��m�SN��d&rܷS:{�%�uq�æ�Zppr�#�&�D��N��G�7���L�{����2P�N����[���f1��5����)@��F=���d�b\4�{~z��޾ ��5__k�|�.qv&mٝ��ç%��}��EG�c/_�$wx�� @��jĵ�>���-k�q��ٕ��C��Ϣ;�I�៍� 6��1�����F��I�����BxArQb�=D���k��*d&>�3���iI��O�P�'�0�$��Jȁkؾ���v�����W<;��썲�}s�
f��g�&v+iYvo��ǂN<*��UpR�_��|�Pu { ߢ`T�����x3XVHÁ�i�E�7�`KBM� ���eS���:�aB���S�";�4���R�(.-]���Y����QV��H����v�c���l#&�"D��:u_wӧ$j��x��F��]3z��X0!%���׻(���y�pd,��c6L�Y��W�H��ǭ),3@��[�N;�|��΂�4L��K��)�;��@�Y�B�x��@��\�+ֻFj+�-�D�u��9霈P� -!�n�U��Bs4�ɻ(��rJWJyЎM0��q��4p|�-x���Fګ�@�G8I��f�tՋ��<���vfHk0Y�����`�GӔ�����=b�W޿��K,+i�BpNo�F��;,ı���)��A\�*!l�9'T�Vm�0&�G�b�L��Z�1��0��<�nСJ|�/b3��`9�i�w$$�vʄ�%��Q��Z�ʑ=�����������PF�X������F�%0>;R'�`w��i�����%�� �X�A���}z�q��9h���f�m��8��� ��Y��^�����۶��ҭ��. �Lμʢ���}Ը����K�W�v�jx�M�^�w�f�o��y�䜖��6ّ����ʻN��I���:��H���Z;�g�s���%�G1q�l�.��oq�%�\9�RF%оY�/źb����S��~�2B�I��Q�ʒ�}hѥ��!��z��t�-��}\��GZK�I�J�f����z�c��W��|��T"��B|����aǅK����T�D����|<�MvF���"��?�W-���#Z�Ԙ�'�^�b�SS��]�e�QL{ks�M���:��1_L���� ]fM��[��a�����j݄6"�f5A�v��}�XA�>�3��	t��bv��BW��Wٺ����<�(�J���l)��%<�}�:M�+�8���nFl]ګ�}	GE�;=-�Ւ]a"�$ޡ��B[�J���$��ot8�_Zz\E'+OQ]N/}ķE��Wcd�-�z>b~�OQ���&��w�x�`�v���<�N;�g��<�q6Q'���/q%����?��3�����Cr?w2]oDHwWQ}��V̥O�����8;j��{�,�8�BK㉬��c�=v�N�f^nS?Id�<��+����$�1�é�2�f�k8�3�^sP8��+�ca��^7���$iB�}�t>@�i/I�!F����{-��F;4��xk�͞O�z<i���֥�_�t`j'@wr�_���*��S�6�6lfW�|��Hj�v��D����V2�J�<���.�"�c	��l��@��/�J'�6�(��!N�SD����k\8�?q�����������bJ�d?��xj����)(AH�i�[�i��k���[�HЦ���,��V�mu/e�!o82�b��'����!'��P��&u�ۂ���Y�W-�%�m��2c��d�����" ��C87�Y<x��N,P�`������q��Ld���*w�!J��m������N�n������>p�.�`�{{���ji�ݚ��D\jF�}7��ᶻ��N�oL�~Uh�u�~r��j[�ެ���d	:aN�%ZjE����6e���~�揹�<i��3�95(Ӝ����z���*B�'�����%Zk��0��
�Ƒ?�
�L��	az;e���}K��Uo�Z���3L��(�{�c�DE�����i��]�NT�`�*|���V�ԝHs��w[�Cr_n Dm�����ϐY�����c���y�R=�q��hl����=�"�WVnAߚ����E���r{�V���+��|s&1���O{&/S�w����p�h�׹�H��2[��*4KF��O��զܨV^�r�|��䱞���#��=����FӬS�i�3Q�m���U+�x�L��jGϡ����N<�NoOɼ*02�����Ok���;�A���mς!Ȥ'�����d\}��b���.���zm1�sQ��2�������\�����������{Z0����t��W8�3]��ӑ�y:����0�S$�F�>���g*(�4�O�p�:h�n�=|���s��ԥW���u���0�h1n��Ι��t_��j�.�u{t�܃��@���&�O�8��]Z�/�N(_����:.0����K�Q\���ߠ.~Ԩ�q�h�L�[��#.�	�^�>0�d
�&�F<�O�f9��ÿ�mJ<0���J���̦������W����SFt,�M~O��Z]�0�G�M�^�T�M-t2�����!���7�0Z�"}��8�D��f�%#��i���肘�$�W�([����Me�
1�m�@���g���<;J+
��~�����r�Ԭ�����A�}'�l�g�鴔*!�wz<�e,Jgʻy�`�!��IvF���BZV9�;u�iD�������9X�p�۷A=J��Fb��r��qG2r�:k�n�9��q���R��W�_J��O;�*&��u���X���K��C�3W{I'�+0�Щ���b|���[��ټgr�e�s�8�wΙ$G��p����<c.D^��J�(��3��12/uw��%�W:���U0�֨��8a�s���J��l�B��.
;詔vX\���/) ��=S?ho�op� ����}������U���E��^�jc�g�yY	�^�/ y�n9r����jL�VJ�ڮ��5z�ڱ�D���)�V'���x?��-��P�>��'���S_��q�>�u�O�&��V�8e8�Bn|^��A���O�Jc�]��.��d�^F���WA�@������1��P
N�N�c�n�t�8��T� ����)�&�0z��tf����}����.GK�o`��� =rW B��@�b����k�ϒEv^7��cȚcɿ�!� ��鬴���1_C�~mi���J41O@<ȸ~�c�\�Hυ�}�#%JT��el�8�F�Ӗ �`NR��S�w�[�\!�kh簎�a,Y�I��Ɂu (蘭�~w}b�J�PN�(�������\:����;�:��o�8sRU�	�R�?os�Dw?̘��E+^�rq��a�:8^�E[���������+<��W�z��2��w/?L�����5��VW���Yt�(��{�7��~�����-Ҽ�籫h}
6"�x������d<�˂�$У�=p�&�B�jd&*ڭ��V�~ -�^m!/8?��aړ�ks�D�Xh��kXf����ُxƷϷ�/#�����0@�+4u?���-&�F�n;zt`m Vb\>�ȶD1}N��P�Qd���V�P��� �:�=��W���=F׏����wOT���E?��z��yj�Q5���48m��3���Ax��1���6ϘY�Z�8fK�u�?4w�D-�`�^�Z0��*��Xغ
6��&�z���su���;��^���� У�4y��Ϻ`Y����<�q	K��A�`޽�������d�[m��PD�!��3�d�ެR��}�~"{Br�����)���&�l0��%�k<I���� O��'&z9��$�<wI],t����ԣ�hJ߷+����/�?����5�2�R��C_x&v��᭩:R�׻h�#"�8+�Ĭl�ӡ�����G��)�O7���⮾ ]�B���O3�y[/*T���͓�ށ]�eЈQ/�u1X��� n�����`3H8']wK��k�ŀ��/��QX����à<ȌD�&����#V��E�=5��L�Z-���>~�x���U����">���@ay����%hp~L�����ط�Jٕ�[�l�Z�Q�3`<(�،����Tx�I�m�����+SԹYn�3`R���v��/�3���몿����&˺ZL�X�C%���Gk7�����AX���bp��P:t�HF}Ⱦ�+�j�z�Q�;�ARR��ҵ\?[�r���sՔ�/�����V���Wt̻XĘ�X���?��"�p�h���K��R��C�^M�� t5~����>��i�l��[~t~��a�b8�*��4���="�gZ4ә�2S�P�<�����xĈ�6��}L70'�*�M�o�����Az�ly	%k�q-`���*��ʿ�F�S�����?��ǁZ��h�!�`�y�}��6��2 ��-�4�	�]�<�h�*�?��.Y�l9���l:�w*�%ϐxK�Mh�eC�|p�I��i���d I��U�G(2�F�0����0ǋ`�inZ|Tه~w�9����Vi��r�أI�9����!���2���>Y�Cd�����9�h�%h:��&�Z���!.x�v���݈�@A��g*�)����A��d���u��%�J�4��FԕQ���`7܋C7�!�A��H�f*����>��K�L�	�ު��O���k�����_�B[u�W���#'�� lM'�������?F��OV�/�q�/���w�Kmu��&��@ŷ���O��u!
�q�������z
�7���i�%��@/\�B�C�9X̋���D�!��|q|(tJ�_X��é�@]5�l���E��gaH��x��m'�uo��S���.�d�$,�N�d�\� ��,�@o}a1�����O��6_����y���36������c�~�hъzh�+�G�W�1~�D�;���-��Xa��(���T/�˝;��r����V9�Fq��>��"%�$�� �Kֳ���Wj2�;���<#{��ʹx��N�o�&��U��$i�>h��t`�0�o�	Ȭ��#�?Y���+�<�qM:ǥ8��4!�	���[���|�d����
��M�8t��k���?�M�:I�.A�Ƒ&ofPN�LX�����#�1T�plPst�!y��S�����v�t#��L���p�b�M�8�qU��AD0k9����:�#Fщ9��{�pzW���+l��}��+ٯ�c�O��+����_]�ȑ�>�?�����s�	�AVt�����862I?�?*�SF�䏧B]"��c�]|��I����֪��Wi�%�?��PZ�5O�1\"�t�������V"�V��G.�FW�2�06�5���S����w��X5��8{��ʂ#�x�wib���y��Э�._�P�f$xY,�3���sm5*3N�3��h,C��	�]	�� ^!F�^������"ΰ�:�W���尙\��$���œ�	���d|�*T?��J��S���q�~T��A,В� þ�=5�&��,G�r���`��7�mz��z�O���u#����"��
��USmf��/��X�^E�8�+�⫊����k�@%�G�8"V��m�3��e���6Չni28,����ܷ�}��^+tO���+�y�̧+��F)-�yh�H2����Z[cU����������̧��w�m}��"�8�Ɖ��S��I�� F�p�cҋ���^Sj%��>�\FE�ñ�����á��.Љdm�n�^q�S��T���;�G7>~��������N��$�?���䀆v�������B���H˯������%��)QS5V���캴��#��3\5c��F.��Aq�u\[q���aнb�5����ѓ��PPʹ0e*���yW��_�_���+Qn�Œ \/���=ޗЕU��Fw�%P9/4�;��'��aSRx�[����cy��b"c�xk���h:��'4����u������
��.y�p�5i�gH�}%&����HF�.O�3�n^N}�ש�C�e�C�fm\G����Zs��Ԕgw��%���#��o&�+T^xB�ݙ0'��2�ғ=H`jxw8B�TIq��'lj!�ڰ��r�+��R�tڟp�piA��M�h�@[�-�u|��h��[X!��ľwD��L�e�Qa�'(÷ɼ�$K�)����k���+�2�R���\�o�OC���f��3��~x`U��9+�;���)�k�&q����·S�ߗ~L���p33QG����l</�h`�;�ϵ���/���DC� ��j���$ï�����An*��R�Ǣ+Y�eq~�4�7x6�-���i��{	K��+F�I��m�F����Q����?rܑm�D��FB��dM�mO�lv�f[�Y�K�HrK�b��]���YdK��U�G[�l3G[d>���|�2��[���%m�Y	��d���M{@F �
�2����""�`&P�{N������<t�kN�x4K��gD[�":Ӊ�R�7���M�̸�¬�}��P�Q�� zۓ��"wT����|
�% Z���5~���@�	ROE�	��dFG��SR�&WG���eQn,%e������-p�1K\�KQ���AHY~q��A�d�ė�?jJ/<Uo�҇�U�ҸN�A_A�6�N�7�B���		[v0�k��`�'������ݮ֐�եQX(�����j��9aTtm�0z��qr���0�5����Y��kw=�׹����m�D�jC��f�]b�<����0��q��8ܠ8�=��ӐvdT���m:�*�C� ��x�@��6��śk���Mz�L}�a�E�I���|"=��{O�O��_�OM����s���@,�z��!p+�|�S���<_��Jܨ�U�v�o�\71�h�Y���-U�UtS%�}���YUZ��FI����v2ß�7r[#)N�`��j�������������T-�N�l4�DA|�>��y�!��Hy{ߴF��P���"	����g�X3N&4��a6-�ӽ�	?.{\�F�g��E������}��Q�?��Y�b�"�v��]���F1�
���B^���
P�*S�D�*���G���q�w��2�rOKF�[H�����S�v<:xO��j*A�;��M�T��Y� �	�mw�U�a����μ� 4�\T$���dp�p޿1��n���4ߌ]R���s�|���n���iC��u��@�c�B
�͌=�ٟ���g�Y��T6P���<�^���
��A|�&gI��M*,$����xk�b��>���\����L>12|#4B����q�=��S�S���T��|�6!~!a�:�7~��̈́�k�>z�+I��F����b���Sl��P�5m�َ,詎�����F��JNy[�L���b�O��
�X��������u��_�E�o\�y.k�u]f�[ِ�	��ܲ�����6r�}3IG�G�fj�7Jh΃��F���?�k!~:��%�Ϟ�e��r���x��+5��Tt4)��2��P�}`�����#���9�D�t�/������7I���!�xm��>�!����/� �L��3C��yYQ������[�V�@-lGDe�׏VEZ-$W&ݳ�#��°�ͿA�h;��v��j��R�/�A�+lK�ʈX�7�0$�_uCJA�x�R|����%��܊�<>\�3w>x��F$K�c���	 ��H�H���q�?�Y�%��8fJyR�F�C����- y�,4�݅��8}3����<����#��`������V4�:缪wr��Y�'��ڵV�sIx;咂;ST�]:y��<B,a���D����ʼ��TW;ĠNΥ�ʉ�eȷ$����;#�=p�����c"�J�j��	�|	? �`�ڷW���� ���L3M��զ\��2�?�la��W��Z���*4�G/����2�����s�� W,�i���a����&I���yd���ֿw�����[5�wU?�o�Zi_j9@���ڱ�8!�$�X��892�w�o�e��W�#��OP�-���j��m�K��MiѐG;K�؁[�}�e��-�e�o�9��~$~��/܂�Z�~�+[�zк3�%2�%��-gv�Mw"�LjAW���M7zN���H�6�U�7Ŷ�ۛ�¼��?U�=v�Ma^������y��~Y��I���G��;񯐲��J _
�ǃz�/���(��U�U<,Gj�؀��d�h�L�LTBt.�c����7�|�c��)�œyh�zS��"�T�3!� �6���N�b伱�Ʀ(&���`�M�4�����v��V�2� �db��	L�Jyq��=��ŀ�M;��#Hc�Կ���!���戎�Ys�]E�NVC+�RA�ׂ̠%6#���q�Pz{�l�m�C3��H��zH������3�!2����M/d/��(��>�(x��n��9E!�+]4�`W)��l��S�G5F:.E�G������Dǝ�g��<x��Fh�1!|ᇅ�O̊�б���M���M�p�X������򖽰Y��C,��gĳ�uӎ����3T,ň-���lZ.�d�P��SǍ���\e4I�Ӻ*���g3JxD[�����/��e���5���k/"l�.f���[���,�|"�`�<�52^�3��v��W���{��K�/���7��_2��(��;�;��k��ԁt�ӳ�%��S������SA���^�3ՔmU@#��b�ߨQ_�e3�a��z`���ƨ>t�����P�H|18(�ĩ=��� ����H+݃5F+od�E�w����Ț7�h;��_���~e��2!RE����]�S��o��M��w�5�^iT�%&��������ɜ�C8_$���%�}�%���?�6�o��c�CG�Ƴ�]�~���ׅj��4�"'1�)��Ϙ[���� ��2?�Σ����;�����,�æǛ�Q�E�F�R���Cx�m��m�Ϳ��(�g�R#!m�0E��{� ���7��?��.7sf}�)U6�U�#p�:o�;�:�g���[��wYoм�𶧾�(���dn�G��8����.td�*�	�� m�Oོ�sdT���+��s#%�ܒM3Ǯa"�3��Ћ��`�t�Y![t����Mj�%?�TexIB�fQ�fIK��� ����zB�hn�2�n���KN���"3}�U'aP�$H��U�Ɩ�	L�vJ���P��)��n�����V�U�F����U*�t���� ��=-m�q����h�AC��}FJݑ�%�q)A�F��'�x!O�ړĵ�O�"Ok��M�UF�r�,4;���є���}#�nr3M 
_m�t 7�������uT���M����r�i ���XP�s�����@����f�N��-����A^��@Q�65�&,�4���0?O���2�v��_;��OƟ�f�u)%!n�1�v���yhx��O�����]�4��s�Q��0���Z�sh����X����,":(0OB�� N�0i�(Vp	4uJWH��X�%�j���_rԌ�q1^E�O��͜�,���UC�5�+�
���j��Ќ@�Ƭ��`	���-�Y#I�oå��J (�G[�6c� �!؛-�`��y��f�4�i�F�X�b�ǖn�*ft���Ծ����j~d�4\�,"e�(��DԜ=�Y�D:�#Vmߒ�uXȱ�
S�(��]��OT� ͉̎��Kh������N��G����XF��I�0[HV� p�%{X����9�}��y]�P�^����e2�� >�#��ŔB�\�����o �����!D��9`�����f�O������Ho�M�k��/{���M&-�w�M�*������g?��l��ϵ<t�͠�
����;"�m�O�X���g,U���<^	�Zsӑ-�w��3����q��)ͼ�q��L�����{�ji. ]fVf�B��4���5/9�uG����G�:�t^�������q$�i&	�=.6g�����h+���)��`[�`@�,U�x�_�(~��o����{�o���H9ؼ��8���)s�D�=6��ek&�`w�Q�3h1�tS��Dm��#����Q=������6񎛐���z�G�L_��AA<!����v��W��$��"�|p��
b+=]X�ۂj��u��4���P�ʟ7șOl�79D(�8�J8����٣�+�1@�*!!����z��T�nu���?�\��gؘD�X�đ
U����������me���#��g&�V��\B�t��+��']��Ndݥ\��~�Z��jk ��$���Z]��u�s&�=zoB0�������n:�vq�`�).�^yIPcN*]͡���uK���n�K��p��q�h�H8�v6g���u�շ���7h�VƠ$%}~bI�dY܊��o���T��\�۫�+�}�!K�����{E2�zb�����#)�q���OX��Վ)��{�-W�0ydJf�X���$}C���t���jf؝�P͑�[i$���*��'�:~6<��;g���n'��B�Bd��u�8Z���~�?2�h�
P ��ޣ�z#�\�>!�N���[�rXb/.�¯�Y�q��Ɨ�Zc��O`���nM� n�C�V) >:9��(����� H��ʳ�
���%�����1TY�F��m�Ҵ��x�>(�WG������b��r��Ƨ�i� �z�n�>�y⛊^����m�sBÓ�s_9��*��iX,CG�P���>Y��ߤ�W�>��K� �?�Gɪ#�i�#�Q�,��]:�yN�Z���2xYp��.��<�l�JƄ�w�BOu�4*��Ϣ���˜ձP΅�!?{��:v�5���u{�K$�ĳ�LZ0���x���o�>���o�X����gx{jy�8?�f�ދ���'�`��d{������_��]Xq2#�`�W�Us�K�~�0}}�м��&��Hx�DNh�e�/��V�V=O�����L����I�M�á#��F`)q���\�e�&yx�5��ʸ݆U~^���i?���~$Ǆ*��I���w>*���l��w��D�߽Jm�`7n�Gj/�wjpYG��ǘ���@��
ye!T��N�!�:�<�V�����"��0�F ��ڝ�\��;qT.#g��/x�m���XX)�K
A�qdV��N'���&��z1��X>�`K���}��S��}�x3�;���ry���-_���	՛pl�*��+�+ef�Lοd��}Mh���b��#9$|�[B҃R!�)��� u!��M���%�=�O���:�i"i�Ljɕ�;k�3��������ʟ�� f~�݅��j��`%�ڱ<n��4m!�Q}�m��JvB4��? �6��<��B S��^D��C��z6���+|�쀪�X�T/�����99�M6�[f�
�a�1���'�T#U5��?d��6�~�wKg�+�(�����X3���A�_�2��*�i�y��䌒.��wI�9�O�!�f;���ךY�o��#O���+T궔�5�y������s5�,�!����d$滊���e.PΙtb��y~�'������$�IS����7�q��c��n4����S�j�F��?@��g���U#H�9��Um|�VCa�_Vt$�������t�Ū�zN	�_N�X(������yNB8�e7(��}FFq0����CL6j�����p��{�Rڡ�	M�k$�ߙ��k�o��$����Ќem�/lWL���/Ψ=���d鶒{��=ڷ'��5�"��5�&�� �ꕻ��@��roI���~��$����-�*���͆���1ds�F|5/;�g�.��B�=�)	����v�v�HF B6�Wo�F�\�-ߩ�����9�h4�����n�� �,���m���2�JbcSJ�9�{돌� �.Ds
F{��������*_�(+��B0i���^ņ�&A�M�_�hx�������8�t��~m�k��ˋ���v\�}�%`s~mJ�t���/��=��l��'V�͡Q�P�|���Omv�Ë����9�i��нrf�+)�lI���t�3h��ҧ���tg�Y*4Q>ЗO�>!�읛����g�n����:k�5���Ya��a,�G�6�1
���ܫ��qS�E� �r��8�YYn���0��£α�e�d�i� �\�:Sd]��LH��WrP�[5J1b���z�0�p4�ˡ)U{�o �$��M�V �g�_�*�����ɧ�c*u�3N��� ӑ�j�hc���DV�0>��0��]hʍ��R=�8g�)D�/�����"[������*���/0}U���5A?Ip�Q��u.��c5��w�|�}li���}�
��}�-O=�ԧ,5�Y��zUVsvѾ|��F�+iz�9�R����@��� ���8$�KG  ڤ֒:Bn��q�m�L�'�Ӱ�HN9&��^��gh�B'�,���@ݙ��ti=��;!�q֮�J�j����\�߬G���=��J�����\�����S��i�h�4�c�?�ٌnL�|���PJd�t��3����*���B�~�WN-$�EJ��M]�͐J�ڀA�ć��[�������=�d���K�Vb?���Cq�(��daDN�����v0���<�Z|0ՎY��FMD�����ڝ�	$�6,��P��
�DJ�kd��k��͙�MLr妔% ������\�}��\�pہ�&1��KJ(ƽ����,���W���ҜL�E��NZ멘vw>�u��ȏ���jutM��.��Y9�S���ڇ�YN�su(�~�4�!�􍤖p����#4n�����K�ќ��m��~'�7�Ov���uB��nhV.�����su��9+�����S��N��h�����-�� �
���Qz���Mw$t�)����͚G���\��18d��JY�k��Ѥ2����%I���x�:ta�e��~t�s��+a~S�f�'��l@9�fHz��-4�p�V�+T���+��Y����e�4�]��ic��� �.G���Z�&�}Z��*��r�z�_[(�A�E���T	Hu\�`�Z*�?�R4��f�6�B�\�I�ġ�J����{��m�bH��Q�ܱ"�=Uk)(k޾�`���i���9�1�휄�V8��F��D��zD��1WаZ�&�\��������~`��6"q�#� �=g�{����A9ע�s��8�5��z����{���I�� �f�����>�lz\��d\�N��r?�⹋J�9P�$�������ҿ��Wc'�7��w�_{\oy�3���ֳ��I��T��NM$���?u.)s4�Һ]�@�~7����2ҋ{vt���<��;A��ӌC;�}Y���� vs4m7�hp��¨־
��s��,�����K�Ě����d��~�0CgˡS�x�K�@@K/�S��}k��<8����������Ca��k(*۹X؈lܺ�D�����w��l#�S�h���Y6�-W������<�c�>��|�O�Q-�Qј,ciD�1�#ZG�q�t�<�4a���^�_ZNO%���}[�<�8��뉥���I��S˯�K��Κe��*#R�����ܚ�յ8(�~��\R��:�OW�t���$=�۽�:ǈjm�R�d����f��R�P�a:#wԳ�[uYo=�wt^�$p���w�^�$l�-�.uVr�5wW��ř��@ ���	*�Nꯢ��Q	�������<rbb<�dLC���m!l�?%�+�����j�i}��z"$����cG-P	��k���B��;.��/7���
�,n���=��sM�ݠӆ6D?�@��Ԁ+���4��Oc9�p��ߠ�iPg������uD�.��;��C|b��bV����"������ ��G[����@e3/�l�����+񾏴k;]gw����h
#a�,���	�yI�4�ah/�.�E�g+��!��r�S�Z�$|T�O	�=
���A���߱]�U1�.��~cR/L�N�<�|
%�,R�3ɓW~ ��aГ��Mw���*�$�"%��f1�l�xι�fT�S\���1��v�4MPɺ�/�d�>�H3d���E�c�$�&9z�o*��?�R�Z˦"�Lg]7�%�uX~��9���5���}����b҉*�G!6�?���=�n:�"����˅�׍�ؐl,�M�s_�}��5��%̒,���
4	�=^��S��;f���CpX�	'��W��!���B<��D�r���	Lcb�Z��[2�a�J��i�U~�ٻ# v�;��.W��{2˺L�ٴe�@'KB6��q$�P�h'KT�����	�3q^��Q��.��� S�Ѓ��_���=��ܳ�N=sn�Q��5s��9{�f��F��Nx��ό�K��~��5޹��b\_Q��bݵUr���_n�5��d�ƙt�P/��"-(��Ă�R�a@�@��kAY���9.���]�O�M�Ld�t�I3��+��d�G�_�;�
��{��k�E9p�W
{Ѓ��]R���!���۾����N�B�|_�/g�w
�.�p�
�P� ꉸcۆP#[��]�!�1_��N�������Q
0�]B��j��p6�*3�swY�=k�!5�ZO���6��yR��2s�h����t95V.}��s��P�$#�	`�/�~g��`_�<l�+�wB�	0�f�st!�r�2Vk��S�@ӗJ��t�a�U��{Y�2�}˭Wpݍ��69�"3���f�U�s:fTP��y�OÝ�c�=��o�wԣ��	ރ�����ů�ւ��o��Cv���u YGR��JewŅ�ּ}����{\ J%S���P� A��d9�0W�sm��h�'���z�>Z�i��Yk�O��ys0\��u7����6lT(�^bv%q�,iU����K�BOԭ��܄��������tz��1����`l�
��f�HFГ��7��mὦ���ϰ��Bf�J���WXm�d�$���b���t�g�.Z��dO�O��vs3 ��C@����74p���ԏ_��_�_�흼S�Q�H����r�bC��P�Շ_&l1���>I&{a��,*��E�9��~YG�?�h����DP�͏}�f'�zI
��	��G3$e	���"yq#����[�p����ؗ�V&�kЙq�]Sj��.� �_z�|Z�������L�%��G+N��~_UoXM�Y,��x�7�q�S#֔�c�i��v㸟7PĊN�آpx�Ҙ���Y����<�76}z<��<�G��	����Q�g��aBh�86��ӽ�X��O�c\�O�	d3��Z�8)��m$���ؖ�W%`_cg�U<;��g����[�!�-���[OZ0OW̱�HJ�[�eRE4��(,V���'P!�wA����|oGJ��<�T�d��-��U�_���K9�� 5;����ڔ丂�1���}0��	��#d=`�61<�|�����'���n7$E���wi�rV�3��G��U��]�nME����P+�_`��O��z5b D���r<Z���b���4����������r�����x�J����9��LmG���ٺk-�X�v5��N�	���Mᣰ�h�6����9M뤉�+�����]H�#^Uc�~� .D��&���KOOB�x�����w�m��vB��(x���g&I����O�P�|���;����b�L���(	�`��%v�1���ͭ��oB7�|Fxi���mQ���ìu9 �m̠�q�U��������4}��s�Y�,�ͷ���tug�(�B�qrb�A�u��1b��+9�3�^*_G��#^c���U�
[a+X2T��$��v��,X����=v�$C~�/sU���˦{j��ʓJ"��\`��3��0α&���d�*�
|�l�=�����ء�䐼��\����C`V��k_(���V��Gk/�z����U����zN�X�c8�R�#~g7H/���կ"eԧ\�yˇΜ�y���H-�;��C���؎�l��v	�D��lI9�������pb�ǳ׸CN����1/<%S��:S�@���}2A:Y�牵{�{
���x�is�9���1Y�ݽ�3F����m95Ow$����~(M�������3����h��œ���&��%�iGP�o�������E��Ƅ������w�V
�r�a���唂|�#���^�R��z���$]����Э�뉪�O?����E�H��Q�#L1�1�����1� h��]�]�?��ϱ��	��A�/����!���Ǽ̄0:D����a��ϙ�������V�ʱ��M�����$>�wx)(Ǒe�B1�� Z�-D� �y$�����/c���䩶ES)��mF�̾�6���眅Nc�'�r�y*wLh}��Ew� ��l�6K�4����.)��Wg6�dy�'<�WGe�X����9�F+�l��2�T������W�)�䅃���i������E�I�����q
_GY�K��Pi��-��'�[2�Z��?F��$=���ܻ`�(�ԏo�?�S��GGg�[��	+#	
��3Xm�3�0��{V����͞�Ę_�5�X��숐�HA�=��S[-f�; ŕ:�a��hQ ��Յ{�'�Nb����i���-�f�+A�/�h^�-&��IHP�l���,@ܾJ�<�t��zj��^~W���#�ا]P�T("�������S���w���r��	�d�I��6*��RӅ8���N�]u��1TImr��@n�dX]� �q���p��� ���+�h5�/Н��e)ȼ�v��S��s�TN1�m~���hH�q5��2�a5"_{ބ034lt�Z
@�fN��5�SCR��ⶁDX�F8�&��;����n���s��z���Qp�vӡ&"KZ���Gc�+�Σ�wJ���-�Rl1��$p������~1A��L�;R��uZB��7�V<���U���SNB�|t,5���-���f�gN����^o���O� �+�c�J���)�t����nB/ϯ��m�g+(2�,[3mtP9�"|��1�Ʊ��CM����G�7��mʪt�?���f����LX��;��K4���_ɪ��w�>�2�i�T=J:�������@ ��6�����?�����VNڲF��d��r��n�ŋ��v��k9]F�<�!���m�ؾ�T��D�v��'yb��{�t�x�8��i�L�Q�c�3d���zk��J�w�ݨ��f�6��5B������u��2@�w2e�Z�0������7P�Y�i�Dַ����*�(� *u���Ĉ@�щAMԣ���QO���{�L)$�����혾�b��'4�I���dQ�T�-.E�Lqa�N �o��^8%3�sK�Ș4��H�,/B�ci��Xᱬ3�����#���qD��/6gg,��b��8�D*�m`9�-���7Lߍ�E���M֐~a�i����w�ogHSXv�I��d���):,�G 0��}�����i�ޏ[j�C&�J�y�;�XQ��J�]�<�> �cL~�d�b��i�&��E��+�I���f���pG��?���6�1�s�/��-�<ܮ�X��As�2����\V����ǅL��ׅ^>��7k_W�̕�m0��qAg�"s�Lp ��e����yDv�j����EB3X_@�^�rΡ�Dpo>����UhIx��l�\��̈́�b~�u����?�V���X<�X����]��US-����dU3S.`j)_��f��>d�{/Y�˓=��d���\�֗,�,��D��:R��}M�u�1s�8/};Gt���ܭ���Y`|(��}��&�=u�}tf�7�C���|��81�E�\e��%<�LPq �yb�{e/��'P-�a�寍[�ޛ{�뤉Y�<������C⸮�m�=v2����$�H�wx')bW4�P�5����}+����ې�9���?�:m��.��R5�<�󠩩uy�NG��yZ~��2�Ϳ�#�\�d �AL�!'��GH�82�{��C�����d��t/�G�.-­��(Xs�d���	���'
�%�g���/(0^n�$��コ�6����L���H��M�ݗ��{C��7[���������J�XH�����l�(�^A5|�p��zxo#��X�#t�"��ΈP���g'�!��+�R��v����e$��v(�`�D~*g����A�a�j�kvpA��R�u���ڕ2�j������fQE?���(,���0��J�q��������EBO[�|�i_unlW�
~,��L���H@^g��MJY�s���E�<�cCc��<���W
�r���w<����j�/	=���x�J�XS!�������f�
�a����F6d ��lp9��\2V
u�Y�Irvg�#�B�t����]�ru[��t�v����/?�Jp����EZ���6�jE�P��$>wq�>��=4]9����5�
*��YXi��j���="$>MOV^�p�ɝm�nK�6�4D�!��K��tra�~/THۈZ��Ul|� ��:��#[|�l�� ����yx���>�`����[����}��AJ��B���	��]ߕ��)�Ӂv�|��4$H��T<w"�d��x�$��'������<�\l<J�^����VD���%���"�g+�#|�(�~�>������593X%��}���
È]T�&�&@��!ua#�� a�5���v�ֺ��S����~���g��w{�����٦1m �l�>Q��D����׌Dk�o:91�T6����p��K;�E�B�]�)~�e�4^*�˶��_�7K�7-��@A<P��0k��
B�r��[�}�}K8l��mW�ݥ�g���u~A��;���ŕ�Z�����m��"�����M6�1��h��''8�����yu��\,��d��m�U���m���9ěX6{�N,�1�^/_^A�§򱾬��R��")ߗ�W�G���kS����H)،P@˹ǘZf��4���"�1�<fq��ެǓZС]\8�$6(8��{��:|��z�,!l����)��L#���fcə�w�0Z���U��b���}(y�hO��8<���G�p�ː&&dK��ލ�8���Z;��M�C�LDJ����5-�e��џ�QI� �_�/�q��Ic��?C߄I�����c&@^�����=&Kz4�5�Ζ�Br$����X���K,�U���+^�2�sƭH{%c�������K�"�/����S�Ѵ��эz/�gB�l~yM��&���J��o��E��a��Q���[im&��I�:l�9G~O�����B����{K'�/�D��^yJ���kx3l�SEEK'$��צہ޹j�'�����8uJX���B�u��x��\�Xh���G�*�b�)�k�c���_`���pm��%:�uR�� �f4���O��Up;qY�"NceaE:����y��Ğw�&b����������#'�7)e����i��QJ�e�j=(
��'[����?�W�i�w�&����'�2��6���iiB���O��j쿘��]�T�Ǆ��L:��=-�(�Y@{_k ���bO\�"� m�l}͊�������Ǧ�z�)�@j�U60Wm*NJ���څ@ԗ�O�@ZZ[� �SN�.�a�\'��'0�ILؘI$Q���P�2S�c;s�I�p|+��x��1��g�e�~_&הĒ����2���7�n2E��2�Hz�hl�J��Q�X4��a�#��X��K�]Zz���
S�cL�_W���mou5z�Y�!� ��8h+{�����RE�4��L]�"�[�P���fvtq !�vP��'GYȫ8�k���_�"�ԗ4��$�g�Rp�M�pI�����Nt:.�9gwh���S��v��m��$3����!Į\�H ��\?�r����vD�J3��x,v��I���Ɲ,�Oـ�0YQ�$O֊]j�(f�b��O��-ޖMoe�	fs���ܖq��P�J��;!��uA�����M-�@|�D��4{��®ȁ��)��H�&_T�4�"u]��ǲw�QE�#T#�@�,`�s<�_S3���5{�6��y�.Z����5T�a���c��@��*
�������Pƞ���d-�$���X�yZ�M-�	���v	Z	D�n�B�s]+���0�
C�bM�fw�W��R�>0���[Q9
�o�e��V��Z�pJ���E��:u�Ey��i{�W�Bs�hM��ГPo�e`�I��*�C�Ũ8�k�$�b�G�Wg;xl��<8s��ʛy�@�\��?�<�xY�z�G]2��o�!�q U�R�Bs��"���;�]`[br��O��{�R���=y���4�J�z��f���=�ѥ��� ��B�L8(FmZ��é~*���+��Q{;pc�u9L�����M��D_)mmu���@�R�q�Y�m���AjXiJ&!X�QeԎv��$s���7ZI���ڊ:��4���X�	{T}��B~�-��:����ٿ���nH���g#"�Q&�[;�BiQ$����k�Ȫ�j�-�.f�.+��Ί�([�+_��G%RŔV��C	�8��Uu1t"�C�7�FE%��7x;`�q#���%��@�7&]�W�+�~
c����]����˳卯D��,}'����j���p�S�`��=��`O������dW�M>i���1���Pz$���2�����n�����%=PrAJ�vO�E�u�!����m�\���?�lb�N(���8T��Q�4���n*/����7�dz�Q��
�}�Y�AZ�R�B������Z�u��{lˇ&��s'$�N-?-�F�����ϼDua����t4�I��>�Q���g����ܔ��N(�:�Q�*,���$|55��ٲp�������>?�V�a}����L�����=h̶�?�yM����mas�!q�"�k��)���PIו��n��FV�S��2F3����YGU��EK���{	�|
�sdo�`�!�/8Wj�zw�����
v<E;r��-�G�CZpV+��i��f	�F��_��% M��\ռ�>�ݘԶ'�,FL��A�Y��:4>��*���Z���M?r�!�����I���5U���k������m��g^�9���
6��搅�{�ܷ�C��B� ���!�>�/��c��<ݴ�p,���0��*Z!���
�zA�>��nN��b����qh�+Cs�2�}�H�%�D��t�����:AzŨ��0�nv&�Ok^$��ȑ����R�S��ٻ� ���*|v}Yq�6Q��a (�g�K��U�A#%c[�����L��:�����>%6��H��&GI�n�7��c��m`ؔ�`Ͳ�����,���b���\NA.	��� � �������rc��%+�G��_K��8,'�
�m�^սG��LS�Y���އ|����.�e�v	ǠV ���tń��R4�@��^�J4V�^/׌d�o�>��	��ز�ZH����
z�=M�Rv��I��i�+��_u�Ԏq^~f�u�S�3�0)���_�[T���=��R,4͠l�$�;Կ˟��XW��XH+Ό8�_%�9r�	�tZ���0P4H�V�ԣ���Y5��ԱZ���!/�S!�\�ݡ�O��P�0G@�|}F;]J�|�f���L��N�����8�ّ�kC�3��憈�;�l�� ´<W!���Mѥq3L�^�L���i4���n 2,7�JXEz�Kea�N�$��ɫ�F7B��Z ���l����tt����jP�������MΡ��G͎n�#:_}sJ��������R?�F�cCF?�N!W���f�kh�D�X��b>�m�;�|y�%���P{�Ny���1�\��	�CXh��`���:�����"�7Q��IY�f�0\��;|���!) <�U. ���]nl�x�"8ȳ�^�W�F�Uh��[��8� ���S���V)�-�΀�F�[\�P��MvH�1�f��sK�GӳT�D�A�=H�sc[�U^����vX��+n�q�Ah�j��P���Q3��!&�C I��r3,2 Z�DK����0�P����+=&|[_#Z�s����i�.W7m���-�ߴ�gԏ��¶2�����9�;Zw����rQ{av-������5�S'��i��6�Q#�;0��Ž���J��|��@��<�R��p�GI�̌_h8�?�s�xb��)K��V2�"��B�& �"�\�!����J�<��#Nu�U��޳���c���� �~4+��Y�}|~ {�$�[�Yg9�6C�xw���C�8����w�e���ߓE�;�V7��ԭ�ܖ��s:��JC7���1\,�vv�~�$ťp'�w�����X��ݛ��#܏`�O�7r-O�~��w�����?#ّX�	���$�)u^�����`�GѳZ\�j
��қ����=(6=�Gy�G%6T�'QޕㅈS��������9���I��S;��`���9P*o��ڬb�� �+�y��NJ��}">�_ƶs�ݷd'z��@����&�{�0'l�5�c�e00��$B(>���i�&�(��HF���d3GV��)�.$���w�&(�)!A��qgM&)�u�|�o��9�����{���k7(���H8�����ȳ��[��tM5�@��ҟ�(��73��L����_���l�Z��t�\��x����C��&�,@>Į��r=ys�����Z�>�zi���D0aq��䈯<cJ`_��Z���p�J~��k�D�l+����]0[�(�9�F-�����[�c�Gx zg�i�t�����_�������?g�do���R���Y�
�S�1P_�|G֋��.63Y
�A��:JϓK$����厞'�p�
f*{�x��Q��H�\&0|�t[��@���kD��[QM�ь:�cI�d~�߼2��0�X�/0�E�+��`�r26Kqٟ=�Q�����f���=9�*���Y &��^;���kJJ��|�۾�I�:"�~��>�_�g���|"���`�=Pw��(��j�M�>H���]P�SĬͨ�}��G�@��¡#@$�L��]s���yJ����ZHZ�+���6��+
3 X��G�|�e$�T�2��s���טL�������e�H9�HO���W�Qzā`���J�Ɉ���[���=bGAn������x�jڝ3���!�{�� ���Ź谱�#�0x�����Σ�pផ��gy�'�1�D$R	�(�$&�I��
���̴���P&ظ'Xc����F�����1f�k�e�W%g��R���*vM��~��ah_O圓��M?CI�t�Jk����dX�Mp�.!A��)\X"k�?T+�J����s���G3��@�BOB�� ?ct�N�r/�Ozv�w�9/�b,��50���<�G� ; �?����f�!��3F�-�"-p�3��`m9�Ȓ��x�&l�=�3ʝ�~)����Ѓb�Qf�yJ���=����mi���9�i������[��{刔X1� ��~��&'Q�!o}lh2p&<�P�0]���b�M�� g��*�I�b'���Wy4^��Jq��%��Y%v�k,�ɢꝴ���]=h�9�=NTف��(���oJ·#0v��+��].���P����˝"���i���r�������W�Uw5[-W��/��Y�
`���mV��a1���6<g���ĺ+1`&A�z
�\�P4֛�"O�*����pף��H��{|E�%[�#�ߤ�G9���d`�'x�E�B,k�<�BX����W1� �Mm(1�Z����p�X����r�|=�z���f�A�v�c�k\�_�>��_=g}�9�ѶQx�u��D��Px��#q
����qtǰ,�7����N~�����BV�qH��81
��1`� ���LS���-Zy���v��;��ȁ���h\���N���K++�}���3ID(.W�,�G�(�:�u��ܥ���R+�^!1���l䪰G\όp�ɨ�
Y��^�Qm){6�/��M8�tѠ34���^�p�5N�BMl�r&�z�aL�nI��6��s�����^&~[�C� �����[�;�没[��Q{��3��*'�ê�~�s�8�K.��XW���X[wD���5FϿ���}���J��	�ux�9�}pk���f�$��w���iоү��ܝ�v�}ma���KP�S�i�Fp�S��6�[�b�ꕒ#�Z��q�!n�m1mP�TpkK׬�Z�>�V�d��	��C�+U�d�@�$@6<���	5���
�����.~�,����=��HهӆsRi�:MC�a��E�&��e��'�%̀����TE�Q�G��g7EkEƌ�zE����|=�aA�;�������U;(�щ�9<
�aN�Y���5͛��Q:�]Y�� �tm��8�âR�)�c�$8��i2&L��g���L��?�L�S8�R��&��;����Ԡi���~�ZŐ� 'n�����y�.R<��r�#K��X��}1q�n�X�=���SO��l��C��C��D����`��ѸϹ�6a^��,6D�^����P�t�?M>�߅��h$�� ֎������Ye)<�e�̑%�N���L����lC�hQ��8�@�<�Mp7�)6x����j+̛������tM�XY��5EiX
~זx A��y��=���1Տ:�Oj
!�'	��˾�7!ƞ�� ptF����-?!䈅�[�_���%y�N��ȧ�B-��<��Q����v����X@�pkD|鼒��/�NRh6yK]�'�S>Tǯնw��AWY�'��h=�O��;�f?�C����e��-�Y���5՚=�k��l��A��6\yZO#�ҫF��q�"�s��q�vܵ�Y���
���W^@=�qB9�{X\�o�G�~���yna�#�\�h�la����jѪ�-�Q�)Q�+�oy��U��ev~R�+�C��x�8M��3*���S����O/e�Ѱ.q�9�� �4�����_���+�����ջ��2�p�h �$Ly�}tb�lc���~����$3.��Wn/�n������A�g(����w�ioP��vΆ#�qO9ǋ�{c��*��G�@z�1�7���QeT:�]����s�p�R 3�`�h�&H�Xn�A{e������p��4����wM���A!��x��ʭ�i���g��������?<���$N��j= �{�
x�H͛�8�mf�]>4�IG������]�J�eF�pF�٫qɊ��+<~�ݬ���"�T�z~�#q�BV���X_g>s���Vm*�'��4`��ǀ����H!8�I?θG
�T�\��l��m�H�
�Q���O�\̨�i�V�|�ȍ/K�Ap�J�L"V�RF�㻐-��PA'k7��"#쯨�\h��٘@�<+)G�Kpa|��җy���L�r	�X�3���f����T|ęʉ8�;)Ӛ�6���o���=�kƴ"���Z����8m'*���;�ʉ~
íZ��7�1�h���_���{)@�:�7�w�c�5�̘��z֤����1�S>0VŅ�a��)���O�!Z��
1
��&,;��/�pJ���;@5�<w��W�� /^m{$&���5DeM�"�bp�V�
�c������	e]�ؽ��	;*l턛-�V_�ˌ]��8l�K�\�9��'ߴ���.f�ٔA�5�x\�XmN��u[�sU���J�-�#7GΣ��`���l)���

V�0�ۋQ�o'��3��A�b$X޿�SHK��4 �󃨐�Eh|r�h�Xw���2T��b=fv��wڈ�H�?�W�ZG��נlG�P�Y6�-�
�`㛁��R��Ws;�TB���ɇ��(P��l�6��"6��:%���b�DGs�y�}�1��3�lfN�Mㄜx/���}ń�iT??���Ps	�A���?������Ψ������)y�87�ēߔO1�(����`�w���#����%y%�4�h����'�lȵu��VS��Bg�y$z�5���+�v�4P�#��G�X3��TmY-6/엠�fkL{
L;��B���?���򽣳��٣�����Ov�'���f�����њ[�h�p�����0m�/C���v�$;�Xq^�ElDP�>{��Ne]IM�+N];}����@�:㬁H���Y0q� �\�Z?��G*�m׈�������*4g�
�/�?G����k����-(#���!�vr�=����_�u7�2dw�.�5�<�&�a�k\8�6��X�#xB�?|>����>��o�K�2���ddo�|qV��f��ȵ�K��!��~l9� ����"��K���@c}�x����4�t���'���.%����������ƝX)��L�陞�c�vT᧗�`ȟ�C�d��8�w��t��o���/_f��p)DOAJ�\#�ɾox�%�*��d�#BT��P�XCu���~-���V-��t�%�9�w����P=J��B�|�a=� �ԕ�ג����Dj���!Ŝ�sr�w|�(� �W�T�"����0���
��'��w�n�y�ڊ�H�`�%Լ�Jwt'����Ѫ/ ����
����b�	v��H�l ��w	=���qB Jt�$e��"
�7NgYC��CM/�\�l{�)�����+((8�'�b�����!��&���)0�-��4/�P#���"ot/�3QtZ����Ar�S�K�D���
Q;i��{E��_F	D��Ia%1�u6i&�o�(�E�A��ė��i)+BtY��w������k�棷�;��u�z�ȼD���g�y��q�K5�N�����T@��h�O;Z����e+W��ݲ�xJ�E�S*���	����=�D<�����T�s�z�b�k��d�'��U4w�G��.P�b��-�T���MY̬�h�"j��!�@�~��J��=Ƥ�bi���}�u�MJ��W�2�_g��X��n���+7�&� ���Iu0&�uz�1ws{7��"�k;qL��.H�2ʹ�UK-ܷ�ܻaU�=�m$�l� �olY��|/K�sǬ"�7wQ1L����d��wW�Xbᄧ�g�v�:���+N�|�p
;�b�e �U�N�fд?��,W�w(�"�fd{�A=T��ŕ���l�;� ��Q@��E(y�����㿰 ԃYf1t�קŅ��a JvB�o����䆸����n�d��4��4[~���0����sz^L]��
��܌�J�Է^��K�3�#ʶ�/�'H����J�αtF:�A�&_{g6���; �a]V���%���?���=��L7}��.�w�Ł�9�f���j>�i��T�E������(s�N��4�.+5��	-5L,����V�����ぴt����U����a��!�Җ<��:�kI�Cpk�E}Ǫ
v9���F_��9�p�����٫��ӷf�Ѯ8�c6�W�8N�t��TJSU�N��}�O'�ǯ�IU���YU�  ��s�T=.��ܗ��o#y�z�HJR��r�[�
�ʬЍ����$���^�?�o�p'~/�F���}�t��TE�Z_`�^�A�8��o �HU�fP�a��C/��ʢLu���dC���[ ���e��2����r���A��+[��pG�݃a�������Nr�ED�VRl�PMX�G�O�	�5�"�v�z����ݑ����[izuˍKg�n�4T�h�/a����x8����~'�Ýz	��;m�?�؎\Ǽ��/c%��~����׸�;���<Ќ�Q�����sCo�m���2�9����Sm:����v\��h��5tޠ?����p�B�(*@��3x��G���V���S¯C響��@q�0�C�,�����O�|�Z��T*������;����
��,�y��d���$���C�=dˎ4Zg�Ƣ2����(��͕��W��jk�-J�Ƹ��@������L��:ZZ���I�k�Kd���a�4+Wj����'�(�	����m,+�����^�D�	��r���22>���ѭ����,8��d��Q�����j��Zȡ�ϐwA��:k`��� G4=���J!��V�|Sa�b���"�fO���F��"f:� ��F���B�3���şX�;Ҿ�|�T���/�/?��*�����5fQ�&�\J��L'��K[{5
B�i��
&o��\;M�ɟ�3,gtWϯgy�O'�Sr&�!��f�_x�6a��Q�A�C�#��2�����	~/4�OM�:��+�.�)}�9đ��"	t6�*�&Iy�^���&w�S7��"ր���e�z�O�ʕ�I��?��uU.ܾ��3E3A���L5XR�'�8L/7&gW9��z��'ղy��o��DƳBK5��;���wr���D�(׊D�q5��}8 |dO��H�ܻ9�ڊ�y���uY��jE�h;�d�\O��D�݋n�3�O�a󉔠z�L��g���*��ίs_a}�LdD����Åg��^+*�^Lˀ@d۲��*x���.xP��(	r�
׿}s�|Xh��Ck&X�����8�5-5�������:��ܱ�9�hζ���p'?�-�K�y3�Xپaq��4��r@����8�E��GDr��G_��"���/�N�()���?y5�MT�ѱ��t�\��u��;Q���C������!%�L���ȑȞQdl�q?��f���eY������	��y�C�a�<���qRkE�&R���� SG2�
���ɜH��*b��B&3y�Z]��oU^q�G(Z�X��_�vy��	(���.զ���VQ�@4!O`������rV%.����&���ie���O868C�6�c�#(��>\�v>���;����a����_���#�TE͍�T)&�R�/��p���;�ۋ2z/�(�wPǱ �|"��!���ZU_@L�Їd;�?5k� p\Y�sA��|�_,��4�	r�9�?U�Z�pz����#7@�v�r�>~����t��?�H
!��T}�y[�L~Hк�p��k_jM�8���r�3��2��}�<6�څ�6��(�2��c�p����S��?��Cs~Ox���2�_*��!z���2_�M��_��{_y�g1e��@��.�G���O}}������Tfז�ޟ�~k��u�Ga��� �"O�{i*發(W��^�Ul��sBF
2MJ������g��[�9`U��;����6���}����=��)��:�	��?�r9��<3�H�~���T�/����Ԉ�"�"T����
a�@��� �Y��q�A�u��z��XbI�.��?ǚQ��P�L]�����a��6Бd�A��SaM]�j m����2x	o�Z�X�C67��t��܅,赘�KbS���MV��3�=#�<�}"0�ʾ���æ��m�=�e����	�E�|R��(~�)�[-{[���/����n�0�����gKa�!埣7�%�Yݜ��*ڹq>C3�l��*��1�u�"�����!C�8�g��R��4�r�=E�9Q�����c�����!;\�^n�ǟ��������	��8���"�q�	Ϟ{OU�2�Y��	t�1L6:�bW�g�Ү!�^�O�x�9��}��:wx���vV�>_�#/o�rUSԟUFk/��F+�c��+�����V�,�g�[��7E����rR{��-5�r�*�,Sv���g�[�J�w�m��H�rq�]oPN+q.� ��j�f齛�	�DxdO(F|���tx�Q7p�oS���ktE�ű}>��o~j�f�������:?�˞�$�xq>��#Ɩ.J<):>7�0_��Đ�F����c��E_	9;��4�ʪ%Ŋl:M\��\�s}?(��� ��i��kzK>���5��3Ԁ��!s���Y�<z5�[
����7��T�Z!G��G����}�s�W{a�F��;�.@�9�x37È"G����K���� ��r�V?���/���wm��Fj0��A[�dl~%�a��f-��?�~�ΰc�3�G���v�@P�!��^���|�6�E.�4x��P0Hy��1]	���֖�/p
�/;D�K�N�gLo�����ewq���o�9��_�d�	liG�:�t�[$�܎L`�WR>�!p���)'	��
�S�H�/ϤTH�1T彥�W��o�X��g�����Q�e����0:/ߎ��c`�X&lf����fۭ�O��m�o���H�ϕ�����s�WF�7��&
�X�D}-�}�3�C�Җ��/�߹�a|�MQW��m�FX�fG���v�X^�YV1A$p�v�q��:�V�7���e��Po�|�C0!~�.�g�2�s���f��������"�7� ԑ�dӔF�QwB���	��,/yRJ��.d�=) ��`�w������[G�k���.�VW�K<�r��p	���3b�����P!K�w֘���Q;ԖW��1u�:�J�8Z�R���Ӻ#[���j��0~Wx������c�O>0]i��Ŗ1�cWm�x�#?հ�?��%�VQ"��Ӡ����{X� ���ӄ��7>0��&��"��c�a�@Ed��c��;��#������ݒ���Z(�����8���_�þ��jf�T=~O�s��0�;�L��Y��ja3ܷ&�A�X�[X4_K2��- �G��|*��dZ
Ĵ4�ř��уڢ�m�M1'�4#�!�f���c��b��g���q~�i�D��gO��a�P�W��S+13�����`�-�z-�h�(s��a:���\dCO;]c���E���&{�Ƌ-�ٳOYy�����x����������8U?�Ġ��ݪ�yi����*?.�@`��&������?�g�m���{�C����	�y2e`ʝ��-��kD���=�S�h ˹�Y��x�`�B,���-w~VtjR�9�2�0]�Y�}�Zo,�Ĕ��DD�j�h�:�c��^���L&�)�� ��J��4�6�Ǻ#�2�C/�s��q{��q-)����_�$^��G�_��	����t�̛F� �=h�m���CEQ�g�u���3]aǹ�03����Mۖ>ƜxP�f) <k��V&JT�g�� �w�"�5����۫�`K_�����uxױ�~'���{l�#o��c�	��fzX�U����q���J��Zr�+���.*��ܨ�D�r�
��_�=�)PZr4E�t��1O���6u�:���=��ML��\��3F�+0
���@n^,ʑ �|0!�i*MO���~{}��c"<#������1�v?�M�GJ������%V�`
������ݦn��$��GZ�	��o�А�%�=8UK9���ᯒ�=�K1�^�v(E��=�	ܝ��K�S�8h�(+u�UJյj/�5�5k[Aq�ͯ.����WI+�	���d��ѐ�)��Z��d�e���k�yB�]�;��w:ٿ��<���;X�Y���6��4�뼤�Yu��D#��e��F1.�z�h�H�Ǚf��ycp�D��767��{vV$�H�_�tW9NΦ��2�C��FT�a6$��Z�p��H�+�bY�˃`�.S��[���GZ�d~-�A�D{6��)'�/�jҔ����ZHs���5��%�;Q����c.�]�e��iX<�I��q�� ߬y .Ȣ5�cFT�mT�����+J��W��fT�Uցuٱ����8�3l|�b*��r���r�a. ���$�֯��)�!o��|S!��h?(�?�Su �mu����z;�!�װ.ʼ�����G�^�f�^y��J�u�s��8��Op�����7�G ��o��#\fy蹀Q�4�4u-��3^������zHU(�|��i�w��j(q¸EH��1��ͤr�A{�ؓ���P}]}A�.<����L����޴$��0�٦'��t�=x�m��۷�&��4 �D���t������ �/PS(C��k�T%t������W[&���/�0130��_�mX<u�.��[L�	W#Κ�ݱ�bjr�q�0��V��7����W'�
��y���z����[Ѷ�*��/p���A\��X>���e/H�G:���^D�,� ��+�P ���1���ܰh��73�w����� �8f4y:u6ew���yT(W��}�����ǝF��.ҷ�1�xj7��9��h�^mh Z�!|�_��c�2������7�wT1�x�h�Mql�v^��i:�{+����:r�}��,̑�kKt�k�w
����������и�3�"���e������o�^�-M�y��y���LH���<�����t�T<!붼!]gT�H�^e��B�d�GH]a��
჌�*	��N�t~��A���/i/���n>\����!rH�|l�(�0��e�(6�3T�y�
�n��`VN),D�)��̇��Un}�H�����.����F89H�0v�v���|/��v83%�Ȣن���^u��M�v��G8�Jbn8�����	����]��9�B��G�P�!g��$BK���s����qgܮ���3,;p�,�����G~���<牔X(�֯�av���LdA�y]c�Ԏ��\>O�hC��Z�ů�b�:0v�d����k�a_��b�E�[��U�oŜ�Hg\��t5��Z�%g�j��u�|�k%�hyR���  ~�p(�fa�T�z�|�Â�e�'
C�tC��6�pK��k�nG�&Q��D�wI�\�W�F����h�%��4��^��I��1e��.�@���Ɯ�ε�o����*f�mv-'P(l{���%������C'�V�g�_�Q]��^6g����qZX�M[N�o����8xS���/���P����_t�Mj�󷌉3�O:]�U0����S�8Gr焕�}{;'���Z����*�M.C�P���Nϐ�c~Ģ�G�m�	��)�;�{d�k�;ۼ��qރ��4X껛�_j[��\�R|}��<�`�π;�˵������
�A5�JmAK�=�H˔�kRNi���Q�{Um=��kXމr�
��n���*�8���L�e0[����`&}2�P�[2�E����ߥ����i[O���~/"8G�m]��@R#	�ր���d��V&��B7����ɖ����KB=�H���	�Pb�*gVT�]D�Tu��[�`����DE���p}N�a����L&�A�yH��{8}ʳC�sZ�]5�eG̖4�5�xKlo3i�\���/�/琳qM2C���E�3�6ޟ���1'�țXw��Vx�bh�c��@4��@�1��k�v�<c�03�$�TIMsV�
��^%����um�� S�]�+-z��e�@��ooC]��2P;s@]�q�_o�-X�~!{`��� 0Ci�Ic��ɀ;��(�*����m�9*�Ʈޣ����Y�Id%� �:���6�Y\��9v�*�<�C�!.�!r}a<�M e���g��
�MX�r!;~_w���<s����c@�V,��ǉ��b�v�6sې�t�%�h�(�']�����n�j��k�8�q�2�8R�(�S��"��O�T�l���=6*��b3�# ���&F\+�O��j j
�Y��u���e`�Z �56�B����(ED4���X���J�d8P���uQX^NVO�i�ż���;Z�>0����"�ۯP���}F&���I����y��
�-#j�Hݢ<z?&h�h|�;RfQPeV|9L��� b�H��2�)�Y<ȃ�#Z�A����ۦ��.�/�!�<�檑�9�ЈV�g�Y�W��.�dC:ٷ���EZt�>⍖��wx�����w![�u�:&'���Tr�j�4�����Z�!$6�%�q809_µ��?�p�}v�_3�TD��󀄫�p�yr1 ���ڢ��K����Tr	�j64t�u<W�F�2�7=�"g���>���6u��ڽ��c��2w��:&�R���j?H���.ﮤ�11�����gt����z8�:ۆ>�Ӝ�>S
!���� �э;���l��~��i����M-�ɍ����*+3�[I��h��"�f/R�Ed���P��X�ET�7E|#��Pc��U1��֎�Ы82n��2Q~M��� W�7�+�n��Q	\%�xF��!��2�^�Y����`�U�:�6	��;5qLΰ
�&�2ډZs�c�0� �B������c�a���芃e^�O��A������V��L��<�r�ڙ�V��z&8o��ڲyA�w���]r��x�lC�nz
�b��@��?}�^���-�TR���3����^�����ؐP;���juZ[%�jmm����Ǯ}�r��<�ߝ����X�)<T��O��u�+�n�:%�v�@D��b�9�941��Y��/JɸQ��ޠ"'��ا��r<䔒��D�C��O�W�%�M��	��)=��%Y)��+���B'a:= ��]ajO�1TX�PNB�Y�L�E�yZy9o#)鼹��w�v��$h�Y��`��KZ^��o+s��
�`>�C�&r!��2��Vw�nS�V���u�#�_(����� N3W��;�^ڥ���p)_�����3_��\:[e���,I��}S�:�(�\�8���R�q=�{eq��!rJC�O&��^VbtBW��ā�d%��|�>v�{y��.�*��K�ĥ�Lcy̪Z������$_.�O�?�Sr���&���l0	��0�P���S��P�q5�b}�t ����`�� �r/�6�w����������K��`۬4�k���r��;��n�X��B��c�D�E$e�m�yìx��\��_���ǉk�y����mٺ�6�up�P}JlQ�'P�=+q�$=!�`>#�g�&Qd����i����3Y�a+D�8A*�c���9�F�$`�*���{?:���S,��g�됪*��Ԩ�^���M޲�#�q��R�4��윌[�d�|��S�?v:������$"�I|��B�ٺ�ϔaD�4�B��Ju��(/,�s�������9		����T���қCX�_g��8Gs�WB�q�2D�!>���yN�|0�H���e��~�u��Jn؂Z�O̎w���P��rZ$.O(��ֆ딸�)�r��	Q&��������U�ն~�P�������g����)va��,ct@JJ~�w�T�wEY��0�w"���!�|�*��
�<[b��=%Cs|'���\G�>�򣋊�B��-V���-Y��#�+�i(\�=M�ӂ���H+�ōC�$��~ �%��塪�l��
HJ� �J�Y�#L/�@C�����P�՝1��������\��@��f�ú�
C����>Z9Q�.��d:l��C{>�O��!��:�G��a8�Nt��0�MƋn@�Wn�U&�k`�Mrl���2^����a)פ���������/�6�����,z�7�<����\�h���.����vVp�!Zsd��]�D�f��rɜ����]  EzؒԠ] ����k�Ӎ�L׾�|&� �-���kiH���GD���Ӄ��V̝o�:okp�*�A�~�N��
i��d�����?�5�����έi�[�ܧi���u����i�碉Ϗ��V[!�v���%��ߌ�Jț�h"������L�wz�(��(j=G{5l��uNŇ?]�l|˻駆ɛ�������$E�|·g��Q�����=��Eǁh�i�c�;Lq�[&��a>Z���H��}����5�/��;{����6o����b��r�V��V�$2h��?�`fCz@�Ϯ� ����FzZ��n @R�5~g:|�zQ�j�����֕�����&�[�mK��*�9�6em��2�'�F��g2���W֎���g!��SM� �/��Ac�"�0SR�4����_�I�<N7�d "K��?o$�#b���x����ݛ"���7K�@7�i�����*��7H����^%�G����_΢\�\UC�Y�T<}�*�$�c���A���+=YF�H�mLn�\��=��VX�0���:qK0"|X��`GX�	�Q��$��E,t����2�?�(���mwO*Ƒ�֏@���X 7ި5��/���um?�Yl�#y�g�!�jO��4nG���V��e*N=P�����%�m��dۉm�Po ���xΏ�ѯQ���=�c29�����0��r6:��5-��8�l�(B�H�E�'�s�9�os>;���ug�[Ш(�0H�oQm�/����
��!�C��ھ���%SIx��NS,�b��?.�"
˩^#dy���ԗ�4,��}6X�p:V$�5KX��s���=VS���y@�
S�����o��ëC,0S�:Vlg9�(�0��Cs`x�R鞱�gYܼ�F2�ebn��b�J�-4�������ƟTE�wͧ'��~����٬��Ŧ�Ug� ��sf��Ɛ�����v���'	���� ��L��?�cI[��b0�<}*D�.�D�d�Dk�g�e��Lk*���X�]�GTm�1bZ	�AlZ���&US��q�dMU�y��딮xc�A�"N��ya���'ʦ����&�}c�!w������,Ix�hk9�u��<j >d�E��M�r�.1�S��6}z�S�C��hT��$$;�4���J'�D��+	������������Y�-�ϲ�L��)��F5}�2؛J�B��7�@8]��L���Lh�xi�r��c+J���f
[���'�P�:5�����8�7�QѰd�����x:���� �V�dT	 ���/�?t:D��Yca��r�[E�{aj���ZDŊҲ�M(�/]� N�
�3Pi�j�y'?3�P�X�X�{>>�#u�6�u�p�Erk�ȏ脈4���/��C�)�8[�v�?��p�O���V�2 3&I���Q�b��g ��ڜ���g#��V�K��?�]�(Ŝ[J�w�ѵ�4�k�_�[hD�TF�ߡ�I]PGH�~e����GT��g��g�*����k[�qPuPa֔^�b��~^Ί�$b����r�$��`ܡ��c?���)�IH�m$��JɈ�+�U~ �8�}L3��(��������NF��.w>�Yy����I�������UsW�G�!�{;7��Wu5���@�=<H�E�<�2�O'���_�ai:'�BM/	X>(��
�w���<�Z.�LI|u�ԇj���B΁6�ȇeHc��cp0?�0�n��/n:y�`�P	[���c]��]g�ۃ��-B_��P�{��[�?*�s�!Nq<䌓��OL�M����%>�p�R3p�w����~nG~�������e�Pά_c���b\@����|?�v�����n@�$�����p����z�2��S���\�oY����r���L�P��������o��������sIm�C�M*������P�(��j&��BI��M	��A�`�)���|Ϯ.e�_.�MWf�]��½t|qj<�
�#�xmH�M|����[�6�=���q�s�Y�F����HLj	{�<��"锾^BD@M70���cT;���ޟ�|��)\�m�M��S�A�������?Xf�
��n��
�� ��)3X�6��:�C�����'��^*,��gL3X-S�毌��_��k�۔��	�B���Z�
%��-�#W��DK��نiX�>�(��ݝ��؃_�y���<���.[����7�������7�X ��wz)|U��W-�E�0�Hc+�}$8�y+�M!���q�����G�3AϹɊܴ�ӊ�?����O�"�e���_�s�ErKw���~ڮ���%{���V��}�o�x���OVmg����A�u���)��V�r�����t��'X�yd\+x�ݯͷ�ҍ&p�)�J!�MŮ�6G4��
UK:|_�3?�F��@��I?� �jv/_!���G#($�P�N]��	����p9�s�F��0��D��鴘Y_G}Á�=ގkS�L3��g�Gh��EV(��d�&|�@�&|Y��2�|�MĩB�,^'4��R���$����C���t�����-���$As�
�g*\�zz�.�?�]� �l��ˮ��\#ң�w�^%������/P{���
`��w�zSwF�욖r�6�7 z(?k��r.�y~��H1\�.s�hf���߳iM�؃�K������8��N�A��f�,����l�SAQ�?l�$n���L��Y!A	��E�:�rf��Px��K5|�5��c˰������B�`�v�'
�m���F�Â��1t��`]�����`,I������T06�ap)����d�<�i�}o��"�� ht^#D�|�Ϥ�&���oZ=@7W����C'�ʅ�{�O��t0&[�֋�2mc)n"���iwIZ��L�������J���k�C4A~)��kў,I�1�����~C}�e��� ��T�1���l���8����ԗ��;��{B�F���0��u�-ܜ"{��s����n�̒��El�8<�e�Pt�T����߅Qz�G�m�(��-����N�� VV�}���7>�A���ʧ�9�܏�ѽ#VU:=z����d$�YD��e��'PiLIZY�ۆ����<�\�4� �Ud��z+� ąl�'j����s#K��F[|��بx�*��I��V� �(�F��)��(͙e|"�$Q4fx�I,�c�����]����L���|���ɾċ2j��)K�EV�-���(�e��u���x�N��-��ӥ��*�_f?s���L��������;���t��M�ɏ֢V��M�JuI2T�s��:�J��;���&�oK/dc;S`��nEh��ځ������R��p"�����a"�nl�K�}�@�"�d}=��.��	�DY���Q� ���
�FT�LF�6�pn8������C}�=���N)��Tgnb�
�np�V��I>ݳ�<�"9��_tԑb�MI=��3�N�74=m2$q~c��*56��ӔA�k�w���9�Ŝ?2C��ꨓ�*���Z�mZx��6�o������y�6�I/B��zy���,��-U�&��֙�������<���`��='��-�n,�ѺZ��(�ƶ*W ����akVC�7-ҍ�����\խ���`;>ґ(��G����o@6�;������ψ̠���������!�1q�c�uD��mw��ӹ硂.�79k;ʔ�����11l��˥���t�ƥ�����0?���v��ߙ9�W"<J�_?n"*�N���.�z"S�|��;}�	�	Ѹ���$���\~&�FJV�?t���u:f+��ө��U
��t^v� &�&��j���:`B��mh���~<�+)O�Ƙ�|�u�$Iz�{���o�co��`�E���*�`�B+��
Y�S��8-��i�H�~M�	j�\7��_�?���O�����M�v��8�p�������8�2�F�[�j(��jM�y�ͬ�,�O�g(��4 �!�˳����z�qO-�%�W
�
H��5_��8ei�,h���A�:�ˀ$��x`�	�?RK�0ƴ��ȋTu�0�ԟ�_�����	����@��w
|�]o:S��9�<T�VB�1e�Qc@fO����{%=|��.3�x[���݌9� O��V����mKo̄j-yw��j	��}�,0T��((�������A��x����5qQ��L�e�,���B�Z��