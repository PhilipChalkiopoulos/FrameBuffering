��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��mX�Պ�$��0�s�zw�
h���4���.}�mA��,�d��e�%:�}�+��H������u����]�jז��S[�"Qc���qiS�kDj`�����7�5G��Ξ@�n���_d� "�!|E\T��C��o웑��hk~A+�V�pt�����]��1W~�DU��C�]|��{KN}����W���ܤ�5.�}D�y�ƭň�a3?��}�g�,z�}W,�ՈC�b�)L��
�S��лa���F�T�e��e��~
�%���p�����I�:�Ң)_5����t�z����5a	L$���Ռ-����#Ac��ŏ�H��ú�?�`�����K/W D��q2(ʜ�;��@���aC���7h0��Ո����D�q�U�Bx�G¨����z���̇�5�/Z ^�S1���dًǑ+����y)`G����"}r��4���v�/��~䮅�ę�����YFQ���q�GQ��zp/�)�1l��9��P���	��KH�����O8�kp^���r����rrȪt��)�I}�#�g4y\�8kg�Ǽ��?�В�;t� ��m��7 
�ܙ�Y�TRa�������^�{c�~_ �FB�;��^�W�RQ�U�J
nL�1ce�8���k�'��Z�Y`��E�=sl���23���Q�F+F�{�S�yIj�+���
Kfk!���Kݩ�w¯Q.��U�^���.M�o�����T���p�h��ow�C��Zh5B#EX(�_���D5� ���Mq�v��ó�xy���K�c�i�]I��%wUU�SB�v��_�9�Y�������K��A�L��H��r���H�b7�	�-��b�o�D�M�/~���u*S&��g�E��U�L*��ht�?�������o���M%U*ewcc����L��2 j������X%�F��nސ�P7�N2z4�&��KG F_���%�?�(������?8#P��;�Y��C!DByDf���{hF�$�a\[)��	;�[�Bķ�Q�m�Ү�����*F�\�|��ew T���i)��b%ڤ�PA$�/�?�Gt]bcRtݰ9����R� m��T� �}kM4wz��4�o�=2|�,�D� R���6��mya�-�	�N@F�a3��ݪ �̬>���RL��_P�m��.�b�b�+���f����䁀��"f:#��6�0���y�ʝ?��4Eb[��<�M��pwP���5�#�W{aM��L*��(�~�H"N�2�BAW!�֌c ٲ�$�	r�IL�"N��㬀���Jk�3�̓�-��K��/W�;.�K� 6��ȍ��x�h�K���T3�aՈ��R�r��n:p:M���6er�e�J΀,QNd���V=�{��4�S6`��[,\��i���p�"��-�2�e!�g��	�3�"e���p>�����˟U��2�9b٤fQ���gT���.��Y@5b�e����M_�-����x�yk������
H<��S]��k[��(Pu��M�Ͼ��&�l�0[9wk<����������J���j��9�H�㪶"$�l	��l��j��
�|�Ux�͜&<-�ox����ϰ(����J�91��(��7���D?d����:pG�_��b��J�1FM��P��YC�	}���6����k��8YL,� R՗�#����š0P�p]��E�ޒ���W^���Q��tNY��lTQE?EE�p���FcfX��#X��Y� �����I����G&�,-2��`Μ�4�:�r��_� �?ev��7�f(j�3�rB�4��3�.��Q�����N�j�Y�E���L����w'����?��?�{�����@��T ����G���y2��Q�t+/rG���4iUZ坸;w�V���\J��&��Ӗ/����L=b������WGǱЌ��0��gq��dq�D�Y:���l�4�'��,��Dw��+�9��-v ����'n0jdr�����j����n9X�>F��} xA3xu�d7\�.+Щ��m[�K��Ƴk���8��%q��O�����N�l���ȹ���AuvB�V�ڋ���9�y����i��7'��$��A�a�3SW淵��!���9����u�ԉH/zmQd��yn�t�5���4������'Le�
�`t�E0��[B�BA��d�����/�D��:T��#�Z�ސh�3�e<2��7ht�����f��Wi�D��t֘�����g��t��p��:�A0�j`�L2�[zt8@
[fx,��ur:����N�x�@�(TQ��+���e��c~��i�����)�%��&N#s3��K�~��łpť ��_�b�^���W���'�1;4&�6:�l,�����@Fշ��Ÿ�p���%�s��gJ^1^�s�OY5��� ���;���/`�x�>Ge���O�e�m��`w���/xo�N���Nh{��K��I\��
�͌�Jwo|�S�8�����1ؒ�gW����Wp��Rź�r
$d�o�ƂfU#��n[��E]�/H�!�Ll�0e��z^��}q{�1�^3m���@w�P���^&�인��&��/E��/�d8p����8?=�Uy�h�Rf�/����B���|�VT\��uK{�l�Ȼ���f��6�m��p�o�J������E�]�L���I���\�Q�a����q	�m=���!�+��*����u@�2>H��b��m�vY�~E�v7~��̠ۢ���ZV�����.CRC_�G��6rj���LyTomFXb�G�\@� �Q���x�`��ά�D����B���+ĎԂ��2�i"t�H�!ҡ�uh�w�V���9c��J���0�y�]�����±�9\c����.���ŨM�c9��T:��N�����J�$�Ԙ�3WWX{�W�˷Ц��s�:�H븑	e������.�^�A�����_�#z� dC�w��O�����ܣ!<2��Mѕ�6Q�
������H��M�����b�G�"��aE͍���A%�$��������p���`M���+�y��ծ���d�GqV�O�s���y��J�Ҙ�l����M�@��=�&_��Ʃ�dq�f�yp���z�i�T,a�^���9�g��5沺���`�erS$_w���&����,�}[Z[9ܹο�7š���8�U@H�O8�o)ݏ��ѺxBIKyh7sL  X�@�L��d��{������5{���^���D[kr�~fA�0 ��+k�a�N%��Z��u��n2�� ���,Uz����t�$j�}f��X>L:�GқZ�⪓���/~��`�ɿ��5��P?e�&Rٗt3��o1��j�xT�}��=k�6�0���Z�x�$�'�'̐��7Ѫ����[�ܑ^�3�C�#{(��]�H*�B0M=}(����m�s�� m��}fb��cyp��Ua�P���;zx�^������k�v��CfG6�y\.�˴�9�^�p�v�mh��sk�E�g�\D��m�PP,�i+�A�;L毥�Ʒ����d`�"�J���n��=���@�����	����H~�/���r=���i�茎 �/�_K�)�swVd����esv�%�W�3W�7U���^��c���f �Q.�r�T�u���+�r�㦈�ێ�B�'��}� :��Ƈ��9U�H�\�_TРK�_ʺ��[{]�p�&�qϾ�����W��B]bx�f�:'>��?��V镎е��.'�I�L܅��KK�G�aZl4��+oD��Xh����1����Sr����O�S�ʟ��W�R,W&�P ��K�W��>�v3�����*�\[�_5d��U@��]?'�}�M6���5F�B]�tM��IA=f"�ؕ }��8�� �N���(�/�߃oP<�h�e(Ob�pv`����-IxI��5�w����ux«*�"��V5�l�c6�>�j��Q��S�и�������BA����Һ�I3G��|h��R��{IT�U������P%m]���q(⸋�$�����d0�G�"� �"P�� E[����u�4Ѣk���R�e��2n��+��zC,����� L�Jb jH�o��SE�������@ͥڻ���}�7�G#���1�"�#�>ƣd	-�{;;��Wf/����"���2&���r��`�,���G�'p�Tn��9���]��@]�Y�TU��A�Q���Q��L.�H!���ꨬ���J���!�S�r���q�3ͳY�'Q�7��h�e�R%�{Q�1ό�Kp���f�?� 0�@�m����P�����aL%��LMT��L`�xX(�+w�K��%���X|��>d��βry9=��M�kѳ׮��j� h�g�	�Gp���;0W��Q��_C�2�C�:�g�l�q��S�i���?+)wg�v�N� U�Ѩ�(�+�l&��r��M�I��P�[zc1z#,i�5��<ݮz��S���#�-,+�,ku�o�i4d�-��I�WF́��M����,啓{ا����
)�]�A�%�1X�o-�)�f)��*$��ȕaˎ?�̲�r�W��w3[�kZs���q�d�gM8ٰB��9)�ӵ�p󞥔[��H=6��b	)'u�L��Xª6�jV U�k�M�ݫ��u21������/���h�1s i�;��7e��~����0��)��u�Q9w�@<�k�p�h��-X|��ϧмpdѴ"�Y,A�t6nrr$A0��@���#|���pШ�G�|�(����FLE���"�s��&�:�N�J/��C�9NQ�����[��\�Q�龞-k����f�e��}������G��d�S�VR�Y_�v�c ��l�#�Mi<l�o,�9��p��䡈�e?�:�콇�s~�ZIt��a�tć�y#��������V���Z9��z&�(��>���E��t�LbKfQ����j���¿`
X������@k�D���=��
(̇*�e��g���x���f.M>z-���ٝ���]�)2p£)4�c]"�RW9$�X����-4�-A<� oQ{'}��Cb����}�j�x4�-��Y2;�0\�G�8]��j����v\�Ó�2�Q��k�&�`>�q��L��&��P��XZ�jj��h��U�ɋ�����	�+�e|_:��X�A�6[h-K
kOc���IY�[�,L��˝�څ?Z͋�%���r��y>_=/��5h������GZ9��+0d�EƼ��6���T��m��j�0~��M�}V�[�@*O����E��J���{B�o�А8:�6qs�,!��yFmʒ�#���֋�]�45?���_3O3���͛��Q�Nyp�����/���$�j<T#T'i�\{Rӛ-����e!f��83�w�O��P-�)'뻋�N+W�KҼDG�4�`�Q԰��i�TU�>k�>	R����*������d�z ��3�	 ����ٛ�;���7�5�.�7ǩE�|d����e'b��b"��oK���Yl}����P����`�x��Ym�zL�40]�J~��TE��;5���4��ՠ#��V`�S�	��а_��橶��c~|f.��!��蠕n&����i�ch�'u�����q_P�cx�ȫ�$7Q�P���i��I*9]��P�t��Q��G�����c�i2�1��u�?�*�Zb�����98d|>��s�� ��N���AkV���GeF����U���/:A՞�o{�_<6�k�ͽ�B!bm)��tȘ_[if�r��xM��D��Z�^�"�1��O`s<ƫ"��3o�3��.�r[�Z:���� ���1��)/ۻ �|�/�10����t���Z<��F�֨	�ֲ`�T�14$��i��h�8��_۬��ΰ�񍟞�S�lM�����q'}�y���~W zaY�-7�^�2�9k��������(��,�k��s9F�Mٍ����"�"���D��r����އS�C6\@e��$�aVI��2��Ț7���c�-�a𬪌����쁖���X5^���I�@��9���1�O�d�G�E꒢�JU��xb#f� ]�_���ô��)��>��rD�����~�i>�{j�����U���Emn�!!j�Z��zFJ޺����r���ѣ��u�dXg0��e��`k��e�_}Z���:gw]ƼUG�s@����`��9m�g� �&[s�#X ��{@�B߉PE�3�[Ra�o��n�0]7�In�m��o���tt��}/��u��4E���CE��ޤo���1;�8�OF�o�q�L�u�Ӧ=`�;�]g��/F��|�����sN�W!	7�"�W�L���1�j1�ߧ�nnO��.GN�Xa+�Ժ&��k��Z�jCC�8�0@�H����g�,��a
:�S�PGy�d>B������+)ݹ�Yh�z0V_�z�;���uu
nz�z $Y�e6�R�?qć�֖t^~����I��Y��q�U� b��zw����R��X�n\K�v �}Da9`�%bњ	�2T��h�Q�6���7��gE,�J;El!O3�Д<�����ͪ[
��?^|A3�e7��}A3�Ox��#��!
�Fm�ejl���L�HI��r$Ů_�\�W ��K�<�o���b���A��6B�To��>Q!Ǜ����$�&pl��)fxf���]ջ�
�k�}�8O!�A5^��h�vI�{�h.���
�$���H�����L�]J�l�y1�����M=�ݞ�l	87k(���2g�D	���$������S�xD&��+p�x"e��F b���}.wG��)���]V���n��p/�ȴә

ϱ WT�=�^ǲ��D=�/;:�6�,��4դ_��]��-[0]��X�s$�����$�3[�H�h�V��-��C������8i�e��χ��Cckxős�m�ed�
�C�^��4���WF��"���O�Q�7��/]�"�����ïU���h�/4yV��$�X�:<�je@ߒT[��@�7$������b��+��c�+?�8JG��
P�x�j��!�h�w�W�t/x���z��=���p��u��·����tqm��Hj�/�8�`^첑����L)@�d�;�S־�L�F/�a��������ԅ���E|�R\@7�b1]8�T'�p��D}�a�X ���]�R��Bʇ2"���L����)���*z6$u�U�Z^!��3��)pK2��(�e���Iv��S��3�w�Ǡ��>��G��� ө��;Q�ʽ�J��u���j�K�I��@�{D� �J�R��d����{�/.��i^vۙ�<1C�gl����ĵ3b��l�ț7L�m��H�a�������|/���[#@g�ǔ�K����^I�.��魖֏�<w��Ё.��,�D(Գ�&��/z���������ڹj�OҜ�#�����u�͈!�'�}��˺ms���9Hǌ!�V�p��f\pg�>E�D��s��R�Ϡ	[�ٕ��s�a�X/D��	^� jc=���ù�4�^����Q�uߪ�.�|I갽ީ�V����Bv��	��TPv��T��Y˟��q�� �m���N�q)�Q�$Ge�\~���W��.Y��-gc)́�LF��B-핕�$;b���P��[���cMD�Y���O\���Y'5�9#�X��1b������)�'�+eE�=���_��^rٶ<������cy�ɥ�%�K�ݚ�p�����_�謗�X����Q:g�~�����O��1��e�v���$A���p�ߥ�5
�A��z`���N����A���}h
_4���S��"�!\}U�Se+�ܘBԓ�{��W�{��
��^����>i>�qr.@�'�bB���ј�����\<���t�*��c�V������?$�5�KQ�=#����,RC,*�|Ru�~�שp"�r���<I��28�ڼ��Ou`�]�Q�j)��>�J��L��JU�^e JBi~Ne�p�Q�H_Ⱥq�<K#����}��c��>o��My5�9�p�Җ��z�H�v1!�_�#܂{Ux ��������'aW���X��Vwv"���萣�2^�]�;z���m�W�r]|��y�(fJ�+��'�O�,��F^\��}c���N_���*�c��9�#ߘ,ռ�]��2���!r�D�roW��+�H^�]?��թ?fK0S��1P�|�*�}�cY@+&�5+��9[lh��LR�Ѩ�(;�p����J�����Ѓ$kDo+�}T�@Ý8���$�8�6G�� T�3t�SƷ��puC�p��E�qГ.�9�-����`}�-b�U,�����fje*_h�R���tّ"��"c����T���"�'T�z�lnǧb�qͮH�;0���)�${����6���4�Ϭ�=�Z�
8nT�I_�D���KST<^���)�
�d�����ޒT���3��g������V���<���sD����wt����հ>��S�tz�`�45� 8�~s���oƽ���u`3�p�9'1�����f�p��[o��p��w�y�w��9���T�(�/s���"�脼��?$�$$ح{����o���3r+��ࡘŐ�WV'Z@K����+#��&髣aPe�f�-wi�Kv�X�X)L�@͐��b���2�@��C2+�6��l�w���y�1!%D���G�B��t������=+�PT{t����+Ҽ$�a�:0p]�6�:��Ǽ���Ƌ(c�J�d�w��!�	R�?��Ys�D�Ht,=`mf����PW�Sk��g���?�h2��QO>�f�{W�.�x���`�U��gB�=W����/q�΁uD�Yl��{2��zG��O5Nf�����C�S�zW!�d�����d�c�<�Ў����\R��1r�:�?h&c_:8*/����V6�d�g�+�RQ��y�UmF���ߦlᖖ�IЕ�+>��S�FO�4��*p��.��E��J�����,�����~���^�+MpXM!5#��-U*P�s��ĳ�f���Q	��X�8�5���p�<g&��,��2����?w��)�-�q}�>M�-�S��r �O|��1W�@QI>�B#��Q�![�Q?a���uKKD�=s��d-.�H�GM��$ҿ�k�ݸl�S*��<J�I��㵛>�2aaÁ����?+ߗ�a�C���W[;����WW��r�!��N�*��.ZBw1���M�kh����Y;on�ɝ7~o�ˈΪ^��Vmѹp�+��h�! �s��XY��5�4$fx���P�d�#�jYË���rK;���R�W�!���btu�� RF5��b0y�`\K��δ��0ya|	�lW60��t>��kO,� �_�I�a�m�c�<�ӹ�ӏ�k&N�'E�������NjGG�TdQ{[Y��:�5�WD���薸{�p$����|�DE�Tü�Ѹ�+p�ʅ����r�]���]��+�{�FJ��"�O���K��4��*&2z<�M��X�������԰�B-��o����/�d-X���s˩�i}�G� �љoo��_`�|mVFST�z|^�T�k=����'�(f,�R6�<8e2��nu��l� (͒Tb�x�~�>��H�/���k7W��[��y��Q�����Ͱ�ֿ6$�0�.�Y�����Du�]��mU z�����f����߲#����YL"���Ϣ^�/y!�(\i��XA�kF,du�V�^���hM�ƥg�����.d���ʯ\���Dn�e+����o��P����0����f�1v�-��Ж:�=(�@g�B�ӝsˉ��&M�JFJ�6��C곗A7���ԂH
%j`�rPd�����CMro������^�J2eЪ��Y��<3�) ]��+�@�U)���ݭ�4�n?�?�Sf���8����BQ��+?�>j��6�ֻ>���ܮzSb��q#�]Hꐮ��Ll�r��es����Av��޻1	�������TrmC��|�������2�j��
�|�����H�v��Ú��ga�� ��V��&Uk����YX���5��t4��^)�,�� �+�ǿ��B�:B��Ro��ҪmO�bf2���6���@qr�D�VU1l����d`�ǅ&��2�<��.�� �B���d�^�����c֮�j�+����� �l���R�x0T΂�����yX\���x�M������P��u�m��ac)at��Ë�ZR�`�J��e�e�Bڎ%v�ݎ�ܯ��c1�8��
���d��۫JVU�u�o5t�<��{=��~�����͟��y	bA��ya�G���/d}4+t`v���/�=Ü�J�y�Jt�7K�p��:�u8Mig�jּ#IJD�35�]�L`����6���Qͩ���q˃qޡW�M<WkBc;�~B�|���(IiBс`�X�, =�n�So4��Ɏ�0�c����s�ʁ�Y���L���L`Y�g����-��yzʫ�ʾB�Xy�w��p�RL�C�z勸f'���ܶ�"�����{)4=���b ���n�p���P���O_��ދ�������mɺSˋ����轢D�C���#t(�Y�jZ{�{q�Yk`ݯ���#WSpQ�S'])��a��g���M�Vd6=6�J���t +_�Kia�u͔I���N��
<�殲�ig�JNj�B�&J�1�Gh(7�BiN��n�^w�̅�uxl�ꘈw���b��[3������qdŒ�R#��L	������!慘1����kS9t��e�2&�Q�- q�����Oԩ�FL� ��.����dYQ(�XZN�x*LT��l��ܗv�}�M�laLgT��mK�F��ӵ�����MlyF�9�j]}<w�瓆R�N:iB�Um�Ѡ�±����ϯexo����E�����5�.�yt�;��T�NZ���wj0�$6��[F(i
��wq_��@pp��F�R�e�'�����V*(�����ID�c��{h+�c
�+"�Cx4K�v �G�L(��g���K�h܌���S���o�z��K0��v��� ��g��f�a9�|�Y¼�c(}-a�U�!�������U�i���	����6�#ç�#}�_ӇL�S-�sR<2��ѱ�&*�M��p���:�i��@^�]Ŷ�� 2߯��ݞ�손����-�������аe�����7�ְd{����*�����Y��ţ�3�����hP�.����o��������?o��.5�Tk[�a����	�M�X�ضą��Aܰ��QvS��y|:��Q\�FnQ�Hhӥ�q��K�	���R 8j�Ep�i�`���Lt���#�F�n1oȄ$�s�ѥL�#wՓ"7ux��g����,�E2'&�Ȕ.��w^D([ԫ���H9�KU���<o3�.Ҥ�q�A����y��Oݰ�ŗ����1�om�D����o}lҔ��%+}����5�o|���o`.��r{��Z��"?�3 ~�K��D)�v�$�PF�]Q��ލ
E�� �9�*|�|n[���\T�Q�(�:����565*7^j�_�H����A����C���Ⱥ���[xWG��ʃ��0�+��"�kB�PB�o?��Fs*�?Ri��ڥ}fl�_5fW[����pF�5�uy��A�+�`^>��to�_�?"Fc�����7�v������e�էC�Pыn,y�t�$�kՉ�ɑ���ݵ�n���n[�J���ƭ���4���]&ձ6j�V�(xXCP�诸n�5�����m�ˡ�:�z�L�G��(���k7߶��0i���k�|�Z���fi�����hu3�C&@vE���p����$D����<q&���~g��z�gE��ջj�;��X�-8�@�9'ְL?�_K���ޞ�H0��ƶ��5'pΛT8����=ُV>�R�NY~��Dك ���y_��A�H7�	�Y�o6��b6�釿&�����(�|;��
EŖ�\��T;W��2�]��\p�㦱��hH�����rŷU�!�L�/�9�ҏ�Qa Cu��j��	˙'d��Vy�>�/=�*yg6�Jr<�*"V��=zU�&XP�~�	����?~W���Y��%V�&YͅRE�{������y�/-znu*���2\��T���
}Σ�|��QӡD\@nj	�����C�Y"�R��~*P{[���	�2���HW�~T�?�2�f�} ��݁�L��6� �FΩH����+��ҘB;�������m�d�j����7	D�"?< �\��>.[>>Rk��Ar�U�{����k������*�RG��GX��jN,t�}Nʞ*r��p��G:
ܻ��it9�r_׶T�7^�򷌇���^�l�O�ӭE����Us�i�@���8���2dN�t["
��t@�E�kz�̀0�+�4�b��h1�һ+)���� ��d��M	�����a��8�Ԅ���CԌ�ZGA~n$܁�*�!��]�����%��-jOa!�-�G�.d�e��~�[�7��pق%q�,��f�M䣭R)����j���J\v�:���
��߿��
�J�[?AO.B�ȕI2@W�Bi���7���(���^(2�B?�~v<) I:T�o��FXר��V��d1���M�뿷,���|#���,7S0-L���Z�e��^4����G��V<����p��ʡ��Ӱ)2d��r��Ws�6�A�g�*�V��U���N��گO9jL��9�f��4�{"�po4;=� ������4w�$�[�k_PD$k̎�/!�5^�*� +p�\|��J.mq�J�B+,��ԓ59�^r��I�F��u[�L�d\x�㖡z����=Qw0F���'{�M��T���]�uާU�)�c��MF��܂�=ع���s�B�i�N���X�|ޭ�v]𝷠K���N������T`�A-�8)���So���dv�T�[9X��0���a��[���x�������um���afI���ya�)w^>�=�gIr�6m�x[T���qg�ml��[X�� ���L�K�އS�)s�P���R�̠/<�~S~�}x�����T�e(k�j1�鈝c�ύ�`V]�"}��B� ���P9�L0S�1�`�aB�Rn2���o�i�Uzr�Є�g�fy5;>$�����٘"=�.�z�_�u�O-��_���-��]%䙗��
�C��/���z
��ˬ4���2�a�V���>P����Α�%l i�<�ѽX��a溷eG�q8�r p5C	#4�ڠ��`
e���J�!��Q��?��r�f��ֻ��i.��gL=��#��O�-n_O10{���ű��r��$%��8v?���1�D�6p�n�`{�ZPPj
[��*qá��W6ȥ<f��.�Y�`=F�Vw�rC6���`��?�$G���|k��RS�?wy
5N���̙/1o�2�n��DB0[5��+nf����������5|3����B�b.HBT�Wɬ̔ޜ�p��{�ڗ��S��{0��5����[�� ��h�}33��<,�M#F��]�%��:}�`�K�egQ�������n.(t�t�ڀ2�`��I�͌,�M̫���O̡R>]�Y.���I���sA�9f1����ݗ��'��{�)�����k��;��<R���E�=ޣ�C�џ�)ݝ(�]�4Vdvr/T��{A�o=��&�WU�f>X�k�� ��ص9�flg;] ����)s�Mq�<� �B��@V߀]��M���a��~x4j�AH�O)ђP��x�Co��K�/�֣OaIk>�	�Z=��&��>N�aF�;c}Ƥ�I=O(��,����]�ua�M)m�LI���Bg1lp����

��C:�����بM��`�1K�:bg�:?W���Q���63�U�1z��r__/k�P(
�fh�Z-s�\�"/�?����a��|۹z#1��]�5+�[MP3���!^?�!E�����B���f�q���wi|��I���,���QH:����<�Cb�'f״�N���=�O$^�����aK�	���:c��V�UQ��ZS�B,d�2� �lO�R����ڔ���#FN�m}_������TM�O~R����ֻ����P�-��qopY���+;����hՈ�f	�ܚā������d@�S��Z�,�.�B�S�:G�dC�{C��6m�>Kf#�6�R��XB Xl�JH�wO<�#fTw����>F)�cn�E�RS�bJ���t4�z�п�@�w��7W�!-C)���؏��r� �8��Y�FT�l�"���"4�+��KՋ9�XLN�����uQ���G2�ԇ��J���o� �J�*z��FvK�>һԹ@����0iW���C�߫�Y�,�H���R�I�PZM[(ŋ=4p�����1|ַ���r" �ϩ��#U��V����"j�(
��,	���)����)R�����˔y��tRKս4
Q�]H��T�ߐ�Kߵ.Z��NOI+A�(�E��j^`�jLөC�(~�lRgG��#�I��w�kG�`9����x{����O���7����"���1���Kꢥ����ι}��;2���$��R���h�|�I�n��ƚ�p꠼�8_��Ӱ7�g�-��m!n�M���U�&.	ߟ�t����P� �Z��Ѿwn��HB�|�1������y�_�n�t�O|�ٱ��J��t�䀪#"�6�YdA�-�y2.��3���a���,�OpR��j̾~l�Ԗ�����&�ND�o���� ��l0�6�ҕ��Z�gFی�iø����hq�As�����x:�fڿl�]�WŨa��>E���Y�QwQ��%m4�ˍ��	�[�@�%:�[@�Yo�U�����U���f�3z%��gh�{l��J���d�P(H�N�h�����:s��}D	����I�<ο�g��bI�NHg��V;cy� 5�=�*C�Z[ƭB8�e��-��;X|5���~c>x��S����4U�{鹛��η�StЂR9>:`s��Q��Q�. ��+P��X��VJE�ҳҺ�S�����m$>�*���ƴ�ґi8Jr�uo�ڬ�&��@M��^3.'	��#U�w6���]���m�8y&�ĺ�%�y/d{IQy���0G]bd�ČȒ�{YFj1�|n�����N�ʰ����R�/�[���#���ep�vÙU�~ѥhϤ�]�֎H�#j��4�)J����'?�#�y�q�/W
��vf�'s8)��acd`W�	,�H����G	�-����/dH���!�%���8��%.����X[�0G�2�g��� 9��(2�@ɾ�/$�T"rF��A��aI9�=$9���w>R���7� ��J(t�Uf��s�-x��D��B�+6���h�9�=���P�k,L�3�׉A������A�Vf��zUh�R�7�B��$�!
]��*^��U'W�B���y˖�F��
ֽ}A
��fLQ.�u�kï�>NK�P�4��;sW�_Z�G�@�i�2;���,�(D0���%S��Xe��{��4�rl����>�Cz���V&�Y�_���%�Hv�����3�# C7+v���;$CF�޹���/�=���^���_0s�u���o����#�ޡו4{+-H*G�њ^q�>������y��h�I������g->37L��M�:��(�u����ir?TeO�B�d}իU;��~�X�s�f��<'���
�7� ��О`s���x�&y�(���.���2�x���YΈ��Ws���&�way���^�ěN��i:�tbQ4'��Uy��ʻW;-Lp�� �������?���M��)r#&P��?���<}b�2����@�s/����w�����`�T��Jȝu�Qcp3ٻ��!�y_!6�^��ڷ"��/, �ptG�R9��]�� ��Y�|�)�h�߰#m��>$9��;��_��y<d�ŭ�Y���g
�FT���ѥ�a��XF��}$�c��rj�V�sj��I&��Mh7�=��wv�y���i����ľP��Yu�m��!�@|�am|��S~�'֍�M�1[�VS�F��pɮVwH:�>�y�W�cD}p�D��J�G �8���[�T�dmu�l��=Nb[��:պ"9�g [n��nMW������MѮ�������N�U=�f|Ni�k��rէyW
λ����c����A!����V�
�ÛؼQ�a�U��#�
��tJ�.�\��^�N��`Qd����5�zu�0-[(?4��b��A��=���-��c����P�恍��_� q+@�K��Aq7*�ca��>~�K7�O[k��rW�3�C�<���d�)����:�]a�dg��R���绕���}� �F��2Y�{G��~B�����&�I J�?鍜)��V��"<m�7w���x=ú���۶�j�/z��>sbvOP�r��i��vO��d����^�ϊ��ڑj��z��R��d�#���C�[������N�� Y���K#@#�ZH����H�c��!k��t������U`�N:e�ɱz�$r	�[�Uϧho�6���|�՝i���[�?�>�6��ڥ��bL�v��1�t u��N��[�������?��f�g�+�F�?&o�1�yRշ*;g��ƒ�	q�[pXg���I9�fڇ����܏Ϟ�~;���V����6�c�U�Q�Tq����U�R� �l���w��x���>cEl8 ڄ�#�k�������y34���0|}����>4h��v}Q��Q���9�`yǖ[�p5k��AW"V [��4��5�cBR@�c3���mO���=5�|���"D��hT��K1�����v
�.Wh����Jݖ���c�{�L����������Am�-� �\+8b��$=V*�7#$}/z�JM���e�"q�Ţq��e����O�ԓ�~'�8����娴Ž��W��%�8����Ԏ�����q��GD�����%d���7[!o�q�rr7��䬅��e<�F��>A��x�E�ʂB5����)9��М��Ȅ5�k�3o�2uH)k*���<j>~��sWS�3���p���)t���	����]�.�;�扔lOw2��H���|f���}%|�ZM����A�߼�Q��-Uf����07���%Ey���s̨�ؠ�Vb���
�[�L^�+n��Y�Zoy.�ELWپխ��H�5%�ڶ��M�g����!Ot����<G{y�k�'�*(W�)oNsc$v��1�H#�I~���P���g6��Ѹ��ƣ�n ��&X��L����{��a���֬�A�0�!a�KV�V��)@z�u�eխ^;'@�Ǒ����_sfPq2�pL8�+����:'�*��Ҧ|����;��w/��p�Q��\�l|��	w��'���0C�j~/��._��`�+���}���A��	��o�oy��_{�+���/�J4��D]"��� �&���RN+��n=�c������uY!� ǐ?2У$�ș���S&q��̌�l�x�; ��$u�5D�8X�*��]�,V�|�4EE����^�J�'�O$T2|��s��A��R�q�jN�/�".�oE/OI^�8���"F�	��D�J��󶛗�Pr����viM���E���?�Ӧù���S������X��`"e���R���Q�K�7��J��˺�ԈX\?�����7g��Qy�͢+ڟ�(@��#M�5p#�E+�h#-�E�Boΐ��2�=�F�][�����$���\>��r�	����HC��D��c���dGa=BI�ӱ o>
ݚ�Fu�-���1O�v��v5��tߎ����P�`���'���7J�_��Q�-%]�O�0���~+�r��{�
d�3��|�s��C�м]�{�iH���i�1E�s�tH�Pd(c�C��Xa���p�#i��)vW	ڷ���%��t�e�8gL�>���ȅ��C��cX'g�R0���M�s�?>.�s57�K}z5�H�6��44�
=���mA���"�g��&}���ܤ���Q�I��c��y��2�n�-��'~ew7x�>�Ł�-H���buq���j`��bH��Ƭ/ٿ�M+t,(��z�^�a�>�S�\�`T����W 3��O���x[ܣ�͒�eJmq�b�~to�_�b���pvO�r$Ĉ2)�-�S	s�-*�|M����3�y����a,`Wht���-(��s%�=�D�2���ܥ2���G��'��ؑ�a��Nv��m��3%&z�_N��kڮD=�l*� �5��N� ��ޚ��"���^`,��{Q�G7UE�?�������91@�IK����ڭrTeU���1�l��M��C����KV����}��)�����~ܳ*��`�Y������it'Vp��� �?3!Z)�����ص��Q��po9e4�J�����2��U�Mδ���<�����4-��C�/��b�`\�\\9��YG���
0(= �w��uV�K,'D�f�/���0��R�z~zoXKe��4-*�_\���K�1��b�د=�^�\I�@�B�V�6_��W>/Z�ɐ�4ƥ���=0��{�3A��Y���b;��v�`��h�G(����J{��ڷ�&M��!���?/,��+�i����/jQ�h��x�՟�"��U�b�����G�
ke�$�BLLF�`7�����+���E��x��ΰ��b�� hlG���V��D���ҥ\����p�3g����',�~��+�V�
�s�����%��8K_i�W&��gL��7��͐��*l}Or�~�S�g��{e���*�	�N�M����� ܤ{@3��æD�e\d���S������ړ�Bi'Sy��Q��x2�q^��+�
��"���Kv�?�Mq7�0F���z��JOD[z{;�5L�_���څ��,���&���J�]"�x��yQ�竧��� �A/ nA�x�ύ��R�q�щM�.�͊`��
�!�C`)�|Z�� l�;cY���;�W*��<���с�7Z���3N%�5�ώ�Y��A0��c� O��Æ�>�f���>m�	�@�Uk{��"{���(�+�ű�
-����Ct�!!��7���=��LR`u �X�f*�}L�Ѽ���_4�f�ҕ�窞2������Z�L!��s�t�Iu������d���9�7߯呞���c���G���],QH R:A�@S T��|�@]��*�Z���z�����j�?�lm�-hM?���'��D����E3�!�o��r�����;�`!(𶳟h�l(1�� 6�g\����P�[
`��������d:���Ǘ��G9����+6Ϊ����g�tg�*=�K3�z�(�q6�����P��4T,�Hlo��OD�TV�A�ܤ����1b �L \8�?~�6
V6�3�=��͐�؈��WS��`��2vp�;(&�5���(��܉i�Q��@7:�V��ڳ	.�����j��L�/�.���6�I��p�-�EL���E��ކ@��@GpDYAg��Ư![�<^]-�`�[��*�b	!U�oAA������7���ֿ 0�P�;޵�c�Yp�3u�c�(/�_����^ď1z.���,�`	.�Ǣ)�L*)�[��{f�_N�[]�(��	ʠ�lT�ix�Z��*�{�WI��Ǎ� #7��<���N_�(�p!���<�T�h��i��ylzf��p��Q*�@ٕ ���%�'=�o�}-P�(\�euB܆�Bu�n�y����aq%�4]ԈMǋm�(���ATU�7b�=�x�߁i�=׷q�W�$ýn�h����Nh�.:��9X������|�e�Qv�@4\�I�n�����Kk{���i��m�����,�5���?|ژܴ!-	�R�����}!Bȣw�
Ԃ��yJ�Fa�36t� ]Z��� �*<bH8��6����r�E��K;��;\[���Y.��'�*���/TB�Ĥ	>��d5`�E�#�L�<R��-BV`��dN���1Z3�!� �x�FYl��O�
\Q*��z�L ��}���:f���az_5�M�'f>y�b�d����L�~0	��v1z�"�!T��_��I� �E
�^Q�*�U�D��	�D�>�]��t,«��'�gТ?i���%��P��`�! ��a�R
e�+ 鎃ʵ{�?E�Y�ۑ�넞�u+㱕����f�XP
������$�1�u��r�z�C
�Υ� ���_t]�(iR
t`�����k|�$(�H �q_���}7��ڹS}S~��c%K^��5IG�'��̥�ƎndW�:��
���������+��NFf>�4g���ږ/�W|rź;�/�w�#�)��-rb��[��֌��;�Pޏ���&)���G6���hJ��E�����@�{�e\�I铑�'j��ɾ�!'�� l�q�Z���H���O-HY��=�2�a5�;���/p����*��'���_�=�����i� b�����P!�~)E�S
ǸbyT`Ve�j���Կ,~�,[�Z�21�/��?��T��JCRe
��T�6J��������E���:;��f��eR���S+�ؿ��T`��'Қ�]�&Ɛ���;�Y��!DV����d�X��2shү�)L�dH�QEF��XM�Ǻ�������Ou~�J��Ո0_�w>�e��J�$�+�⭞�y�:B+��K9{�M}z�\��l�W �C��&��E��PkA	�@����.�[� �87-�!�#����K�Y�+֢-�d��Q�f6NvMB|�$�Z͌�+q8�<��M��L�����5���7ު91�QGH�9誐���󧜤  �v�:�^��.���+y2�R�x\�<���+$-yf�0�F�(��ňw�wg܏AL`ƛ����)���w�B��Z>(����:[L�������'�X�IHM˷�HJHЯOl��=�D�"q̻F���
,y�Ɵ ��E�4*l�Oy�sD,�"99�c��4ňCr��P�!Q�h��u{��<��j���(:��<�jL�� �>�-uiXxO��}7�x�2�7��RΡ���N�Y�9{�x)��ƻ��K`Xn1�u�Hx�`��(�m��D�y�կ������L�}$v���Po��MhF!;z��;� L��-W������\
�(5��׆v���5-!$��˴��.�讻�D�O�DE2�=# PsƆK�r�n�q�r��5�c1O� �*v:}#f�%�?��	ERňV}b��L� #���B���Ũ.R�.&j�*թ4i
<'4�5�t��S���Yn����_^t���=��t=���M7�2����W��r>�&:l����~�����|B�(I����)|��W4��z��`�&�,	�������EZ�g�tq��H�/��gUd2ب��ycHz�������a�g&Ϣڑ�����r��v+O?��ϛ?)�d�3L��ׅ?���Y�Q*�&�n�y�/��U���Ҡ��a3��c���ν����G�>�a?S�v ��C���@P��0Xn��xa�gZF2�yX��}3e�dl���Oc��s�k�O¥9�m@D�f�j�2Je�'�݃y��{7��'<�c�����k���y{TW�0R�6���8�-͑b3��{ �$hk�{cA��g*�1�8�(���Bh�0���S
u��1�$b0��xJ�]_o�F	��s��H+:x�妔��59��F2/>Y�0�2C#nQ%D~��5�l��VU����5�Ǳ�4�������<��ˁ���2������s��U0�Β��$�NK�@�`�lP1��(��w��V��~:��ڳ8^���&�O:��	�F|��I��<���ܵ/���G4T�]}G�*9~�w������/�*�`�x�&���LG�w���y�
Z?Ǘ��=˺�*��$��Odk\��&����[QQt��c�r��'����c5��޽o�|���&�|E2F�ɯ����I]a��O����W��Ȋ-d�O3�ϟ��O��p��I�0|�lGb;[�?^�>����P�K���ӇԷ�،�"���}erW�P�%?v��z��fφ
5�l��I�ض���d8�
0g-����񄢰S+��Q-ڠ��T��jwШ��
�ܷ��]2���O[����@���� kҎ�Fa�ǖz�d�J�P��@�P{�ȏ�a�=ySC��>����0iE@)�$��6���Z�����j'�偆���h������c�k�0:��K^2�`�!US�ŷv�#!EUɩ��T:����2��G�x�/�~�����A���i�#�э_�b%[AK�YVc��oE��i�����(0|�������1iҺnX�\��=�v%�h��/��00����̽B12�eQ�̩t�ɲ���E:�Z�E�C���L.e0 �+�`ե�A��@F�"������<�c׳�7��:G~l��Ͳ�hK�5���D�k���;����]��*�K|�����D&Z%)�����̓!�Џ�|JcqL�>�d���uZ�C 1�R�x��vb�o��o ۋ���E�BW��S��/@��pԚ����v��Z�~���=ד0?���ks������AaI�D��ު��H�{/)`�_n���-������+�k΍�rs ���SS1�Dފ�:�B�}5e�{1��
uH�ǥ�+���j*����'KPG�)�׬ɑ����l�2��t�L��><PǺ����&q�m4����4���?�����>�мU������Odw�B?X0�b���\p��i!o��l�pP? ����?���������9#��fr�xp�����'e�q�䓭j�a'�j��Q�aڏ�ؑ�QqaV�Y������ ��B۸��ށ"�&�F�u�:�����Bh�>}TM�1�#�?��|=��~�$P���)�"��Y��{��E�{��̹#�I�����d�L	�Y���s�v ������Ffl�� A�vb-9U�� V�BN\��v	�?e�T��{�jI�PXk�Ӷv���1��X]�J�f(�Ia�"�"90Q�<P�nF�)^`����y��''�X�
$0��؝��"-T��Z��q��W���4�(��
�&*�q`^̰�x���⟈Rt��,Z��oU���T�Ӛ�z��fe�o3���AN*�5�����ё}��;S�����V�Ft��v�B�k��h%٘�D3 ����{�b�"ӂ?|,�K�LCFv�w��-_�`?��/V�Yۊ��k.�S�b3��4X�/�8k���� �&Q�ڰ�������H4R�h��Ġ����h�{&?�b%ô=*$�x}���&5�����GHA���_�:��g�_+��o�KMМ@�xҧ�lɱe�:�t�F�gz����W�a�	���9yX�ZP���I�Zd�8�c�r���"Q)�	���z۽.P��0x��"��"�I��Y�~��3$���>{k������d������r�C�J�b�o$q9*�7��x:7��`��;��uc��9�����o$�ۀ�h�߹l�eς�_䷽پ��kb9��;:�|�O��� ��Ig��2uDQ��5X�G`G�.�c��Kl _�m%�Do2|dE���1�وwk�9�T���"��$p^���^�"B��d�b=!?A�A��(�r���&�ќdBΪP#7p|y>�*��.�0��yU*3��A-ǅ�h� ����?W,�Fe��j�ym�a��FIWҒZ�`�Z��*��,�dLD��a��}~P�މ|!�$3�.�X��|�WzH(G���7��7���d�=lx���s&9}��I�A1��ޘ�ɖ����q�?nu�[!{��D��[�޳�������=�
���ˌ��`�ʢ��"�?��6�����'��q������Wzf�8�ݯ��f��	n�����j��jj�c*���l��å�m���ו�L�Aq@������m3(q~?�8��Mo�l�FK�.rN˒���AnІ+�[Ύ���>e����c��1?�s�Z�������Kg�}^�$%�W4�k�1`�v-��`��8�p`M�e�O�uô}M�v���)����׿fۉ%-]Z�R�8y�����#O'c��pE�¿'��M�[ǘ$��I!�W'�m�)�)�!kM��P}��yZ� Z������9�̘��_��&9��%Ai�q$������,)\��+1����C/6G�I�J��pt�@�_mr|1�H'�ly�}<#��R��I�[BU��%��a��OF�?�r8�c�p7���8� �隅�fْ���<�k�ьe�ŀ�I>�[�Z��&�O�f� V�L;��*G�}��^�$�xA�P������ݔC��r8����-w�N]tF
�=`����m鱩�n�3��Ct.��w2Ӊ"��X�	��P|�M��3�=�%N�P�iA;q&zϛC��ƪDr�-Nr'�R@0ꉁ���i�5yH���k�U�dT������Н���uX����]D���\�s�~���$��P�����C�KŖ e�g�Bt�M��'����J��H�u��Ӊ�%?�y�*x�Y��;�T�8]M�d4"(Kw�w�R��?��-i��^[�7���Y�^E�8�Y�G�Oy�>K�Ը�N��yz��|�ː�c�909!����9�8\udcUmy��gk�Aa�vhpe��j݄���i_p6�-��o61^�)�?��z�7����9��{�ڪ�>�j�E}lo���@b<�I�F���/0\p�Ѥ�3+[d�٦=���g��WW6+M����&͜k����D����{�J.vQ�
}�ֿ����g[���Ev�ܖJn��"r(��q[l�"�e���(e�b�p����Q Ar��G�:0����7٦��=�B+�Mp!�@ɜ�hR���"N�w�8���]�Ą�v�}}|X!�<����,j�ҏX�Ԟ-�Bm�����
% /\�J|�3�D�p�[� �)��)#��hu��³31Df̮lD����PRŝeЈ��%ؗ������=k���Y��U�E��4�a(8�o';��X2�2�W�[r�46��F�d~�Ȏ3��C{�߱��ü�Td\���S�P��3Lu������F=!�����^�S�=t������A��H�@9��
��a�� ��4qaM�fΑBhWQIx,��FV����, '�trD�7�]T������,�-�p�Α����N������_�� �T ���m�%-׎0���I��$T�������
���M"6�f��ӭ�z2���d#Xӡ��-����OwޘL�Ü�U���<��О��Y�ht�Ht�����2T`��#>oz,���
�M����aG!��ӟ�jru����k>E �����J�L��AE0>Q���?+d� �^�D�	�oM�u�.KHy9'�	�s��?0�K Ow��{���` K��r+��3���0~�� ek̔$'x�˩)N�Å0^^�j��?#t^�@qn�6c�Nh���B[���A�g���6,�4���ݎai|����LQ2e������H�1xet?�eU�f�]�	���q(u�y,>�N6zOÉ��}��m��$^d��6�±OZ��ڀws|0F�DH�#�"������D��F�᠘l��r�u'����L��cy����*P�_( �Bd�I�#8WhrOI��~Z�����x2�i�r�M���]\���ep��o�#c������:z�pSdil��)��-O����{��ȼ~I������+�v;�i8���x�e�|Alg�]W� ��x�-�K�����͂��/�*���<�����[��s�iC��Ϡ2�w�" %^�TS���hNٌ��C��^'g���o}Ņ_d��0��w�x�43�ڷbs-#��LņU'����Sn1APqTGEٓ�d_'(���>����7������<��8��h.����v,��icFX~�m {��1��d�߈t,3�SApje>B��s��E�ڟ����	dan����/��	)w�s8�YǷw�:ˀ�b���u@��1�%a�j��H�ydV���Grr��H��m&�&�`��(ϓCK�ߐ*�z.&�& {Φ(���0�
F���Tl��*��_��_��j��.B����P�Լ�F�`����&s՞���S�}�lw~9���-���R[�f�ߧrS���xo�=��A��֪	(R`�T���<��t)��`>�<O�%t3��!0Y)��|\9�Fl�
;]�=#��3��}:���VPsP�'5�ϙ�~��}�~N��N�Vh#���������p�S���������߾݂F��ƴ{`V�!	B��FLf�8qm~58�*�W�O�d�@��0��B&=x��0���t����f�%zE\^���!3�B��Lu�\a���*B|�Y>@`^�R����C<�ఈU�+�@�`rH��-Q�1�v��"5��Rw*�>}�J2W��uF{c�u~E!pk=�n��8�U�rQ�<�s��?ò�5��$m醅�X��A���d0��5(�m�>��a��(��)q�4ӿ(%�?q`�� NW�-~u�D ��k�C6̘��>�C�C�	"5��ͮv|2�3󟙹V�P;U��p4�۫�i�KP򧪀z��N7+k�QY�d;�����T�雪6�U{/� CHhe� ���R���2�l\�~���,"��j�~R*��0�u�W�ӠcBjčqň�h[���mM��ߌ���C��S�[�iq.������~�W� �<�N؂5R<
��Ȣ���=r��Ҏ����g����<��?w�����������=�
ɱ�� �P���p�|3�Dۍ�y��R��D�C�H�Y����w�C�(g>��ea�n�C�' Z%��x�xX��F�[Ξ�t�Lh�v�����#���Ot���vot�Spg/��",e�.V��d��8j�hۏ@����6�AH�lg���X4�8�n�axL�SM��P�s� �CN�_)ӰQ#f:��� ؘ����-G�u]�1����ʌFw��(2�7vZ.���?88!,u�=~����v6�+G�pZ`:��Y�z��Iy��ߵx;5�^>c��_>��s��� w�ܬM$�v��X�#��Gulh��J�v��M�h>�p�\bt,�o�K�S�}�@�$�h���^�o}�Ϳ��؝�{k�g<tf�o��Ї7ScBGHuC�����iVz&d �UQH��:a�\ָ>�񳪭�'�A����F��ٍK9�r<H�?8(�����Ӊ��3څڅ�^G3j����+�� ��qx*k_4�U�e��{�}:���S�6��΁i=��*X�T�lۃ��$9��\F��%n����˖��7���8d~���ݏ*sw�`�	�������wD\�j��S9+;
�U�d%��k�]l�Ѽ%�� m0<��F���3��_L�����(���H�Jd�]*Ǎy��Ѐ@�S�am7�w�����%6_��P�� ?t͡�ʺ�ˈme{É;$��X����ȣ�^�[s� FʂI�p|إ��,�W��& P��tZ���%�����A�몚2��cvG�:8��"��M_����8�@��ˊ�Z�fg�(m�H$/[gQ�J���3�@a|R!#��Dwڽ&�r���>���L���zʨuE��a|M5H��`2�hN�Y̟�(l�5��׆*sn&q73��7��e����t�_i`#�t��i&�.^f�me|�}y������������C�}�W�Cg�����&T�tǕ�kS�,��B���Wh�2
�"����L��ě~�daJ0��z�(]�`���y�^�n��YG)�쏸�� Hd��q�}Zg�
l�����m��D��vo_YT}�b��w�+0EmR��_��AZA���ft�)|�ֈ
���9���2 x��S&z9G�s>n��5�ظ�V�F�K�wM�6�5�t�2>�����!$�����xl�>W 5��8Ͳ]%��@XQ��5C4擨��jZ�V�h��t�9���*��މ���bF�sa�!�����:�sVrZ[j��lb-$]e<gc���_��H"�爛�{{��eK��?�	3�ܩ�T���8�|�!��l�ƿ 1�ߌ��l��ooN�a�,�n��.��������aY���vj�g}�p���n����_�NO�-�ST�`	'}��tS�aYJj��\�r��6��,]�F��1ZoT�I���</?DqX@���L����REC��HD}���ת ��m�{��k�>Xtۏg�ՍŒהj��f����~��aRF����4C)�u(i�U6=�����ta_`�
��]7'y���v`������0W�f����a� ����l9#��"�$a���O"4)Q�O9}�Y�#|:�*�͏.NlО��rz0����<�Q�nm�n�߾�����sn���l-
A�'΅#x�����z�_}���𔽺WO�!��Lކ�FՏ�>�<�L}e��h��8��6��॒�x��R�!�8�<��ft*R���g��?%��!�(EC����f�.&s(��QI�XxW��#�3i�O��kJؒ��FYL������]�}�F�++���'E����>n���뮾��5~�,����Vf­BϽP	"��eFJ�//�%�׀rm��x��	MH���Ŗ:,ʼU�x�hj���"	���������x'��4�צjCb۳�X^�3,��
��f�ȗ��|u�ڪu�uBH?���N$l��2����W���
�i�=B��P�P���� 3�ԣ�[��Fy5`�����[br̽{�Y�L�o�=`��
����4��cW��ל]��-g��#�7ݻ��f�L��A���b&c�U�<_�6��dϟ�ZzX'��k�������9N�r�1?�M#D�p����&8�����}Κ�(��|�U���*,��;`��en�p�P��T�.pS�dv����~קH��&}3�4m[%�*W(���pఠz8�<���J��K��Ej�͝ W&�uQN��րs�\�s�|�X3�n�RQ�oD��J��[!�e�O��ca8���C�Cқra�h�\�: Z�#�D��Ј�N��X�cy��[��Ύdf�1�d�t�:�VE�xW஑CZ��B�4#M�+]?�iC�UdX�oAu���Wo����ރ����됊r�ϩU_��%Y)�X�K+�q:]��q+効�����Q:ҫ�~���=Ԍ�>�z4�Yڰ/�W'�JJ@����4�G��?�zѣ���K��QG�,DZ��7����`E����_�C�12**�=����˚[���dľ"᥾,�E�6��bG�����]OH�D&>订<6�^>K��~ci��a�¦�`-���6����� ̚�%�e���̾���Q���T�������7Q�̠��P֓w���r9!N���Q�	��kt��P�dQ��	x[��׊��J����ˉ)�-r��?�<mq��	{�GI�#J�#gsrj�h��̀�/p��F\�|�E��Ȟ�aE����.�&��\��u't1�u�3[�W8�
1 ���z�}0�3BYx4��(��x�:H@j����lv��n�c�m�TB�Y��ߔ��u������gnn>$�M�<��gi�{��	���KD76�͛\��yK�j�D�".��hS��@��X�A�Ł�)��߆�!�&C�������(�A/n�'%����p>�R!=**�8(��0YG����8��!�:h�h�+�	+Slf��9H>�|J��/��Hc�X����^e ƕ�z�]�5�8v*��n�3�;�3�B<s�Y�7O� +�-.��v)��Á�H, �tQ�{%zyP=��'`�ks�^���WET\�N�_�&gp��mF�����]������7�џk�	Ȗȕ����wbE���Bz����u*��l�[�ʃ2��wE��CL�@)��$����$M]��@��H/���6���@���O����VA����ĳ��F�tyJ����� ^|	�I��O`�\D�@���N%�%i�b�j��R�c>�ǥ���1K�0`:��+e���T����>��`c�I]�h�<7k�8�Cdr�Ɠ́!�zM�w�(��O�L��)���X1�g�8�*��:�w�u�ӵg�e�3w�����2g���hT�|�7�S଴C���ޭ|
Q����M�?��`y��̑ڜej��Mb�4�q�W>��X�K�g��$g����:�>��|��0������;T�n�k�����->\IY����hW��Q��-3U��~�b1�l�n�!+j��7��� �i�f��[0z�R�e}�!&]�*����=�D��pc�:%��h?u����e����L�
�����S��.A��~�{^��BJM�y!�Se��y�xsy�����v��V��I��Oa��F��;Δ�ۏ�aE��m�n×ς��X����4 ��i�o��e)�)hȘ���{�As	�	�?$�(k?~��xT҃�&�=�Zp�.�P�YV��S��ь!"�I~�#M��9���������a�;�Y�+��z/�����u�x	\b,�_�p| x<���
���.�����L��ʜ��3�ʘ�|`�����C?8#>=�_���f�5uBRJ�^4=8�?�4�DVs8.yH�Z�I�E�|zr
�Y���E��-��_Z���c�(�T�S/,O�:��]��G�Ґȓ�H��sǙJX��:v���$,���i҆"<Q����N�9���	���f���6:�P]�-﹌% �j���f4�j�_j��4����?YJ�fl��g�MI�A����L�E��.��B��b�� �����6�`��a?���dµ4*Դ��lP�%{��1���#�qF�@0Iԣ$�}[M��K'�_|���׻�'hҐ;�����ˉ[��*p����[�vb[�B�]-T��OH�u�"7���w�=���,o�$��`�|
��Q����/�E&t���bt�d aWo:Ԗ���6G��"��o��y���2nY<4%���O�2�MY��1s�'�^���!�-3�B�ULs	_mfi���y��էKSurC
����nn�5�py녷AYsw^'�cV`�����>�)Z�|Wӏ/�p��Mb4�����G�ؘ��I�c���iX�b& -��SA\���Љw�]��΂�֭���t����P�S�;&�bo�׬��1(�cj9�U��L�'���}ZN�������	j���h�%`
���P�2�h��,�!�-�K45��,�$8
=��&�"������ O/Bk��D%��g���� }�xh�Q ��yh�Λ5<��½8�Z�COdӟ�uk�x��C^f�0� �^z�ک�X��a4Bu��F�~)I����8�1�}�k?K�����(�|dbg��#`d�o{R���1�d
$�~Z@DǕ�~�9����qH	捜�Q��[.&%m)[.�2��6u�[�j��F���-�j#srHou%�JB�:	���-�6�@^K�6և��D��Y�5{��J,6��T)�`������"�	_>�H� "�-X����[����m�(���۷M�|]LR�O�t��J��X��X�$�Y��'��B@w����@�J�Q�pZ�3�L��UAEQp����ԓ�]�uVa,��wH��{�F9nnh�ʷ�Y ���a��~���@K
���ҸCbl�ɥ5!NMtP�ť��2�"�F�s�D��%�G�.��>Bio�*<��ca\5cO�E����$v:�f��F����=�Q)�>��RQ� �8�ضi039>��B ��Ѿ��ce����;C>�,����c!1>Q�M�]�ŭ��J�Bi���$�Y�}6����qi����{j7��Y/F�ق
���>����p�Y�����:�C�n�\�9�����4�Yn&������I�՝�ZG�P:���l��v����� �:"a�dG���7��������m=� N�u|jE?v{�|�Q�%�vd��Q��iE�[T8�(n���z���sMZSI^*�²��u/�/!	e$&�U� �"�y`�a��~dFS�=8��R���Y������\v*������Ra����#���2U��� %�%��a�2�rǆ��U-�P���P�{S�M)����J|�5|?#��2|���'4t���	Hi"�-b��l,�P��ԇ�!-ŷ� ���O����V��n�D;z��1�s������;n�NHI��c��G�;qS��B�e��y���m���{�b�(���,"ML]�+v�סA���������1���$ap�B���w��r+�V��{�V�9(}"�� ���/��D9@��a+��`���"���$H�f�`I��g�bԏؽH�^�Ł��:�)���I�p�`Y�c������qA ��Y��
D�`�2q���d���(�D�����-�>~�T �5! �؎Ԁo ~��'��y⣐�

Ys��`�,R���,���4�@��+��(�w\��s��I�栅L�1��W��
i6����M��b���)OK#�׆>DWv��țd>ԟ]�Ы�1 W6YPW8����e�hCF��,(���s����Nm��{�u�p���u(X����s����UE��(ZoUb��,��S��λ�*��?��l?��K[�_u��A������tvb�I��c�	z���K8�tu����_�$k͸C�Za��P� _�\@r�\���>����\[^���4�r��W˱z�"��j֧�0Q{�KijM���;�I:��Z�P�T��Hr�[���\7��7D
�D�E�Ϧ[r��Umf�z�0����=��Kf����!1˦,��W'3�K�!�0QP>Vk��=��k�P���V�d;Qr��D�q,Y������	��ۣ�3�����~���ﾏ�
J�+�ݜ����|�q����Y���I�`�6�����.Ԟf
�wmϲ���a����q�f.��Z��M�\����<���t��mB�KT*�Y����މ��6Q��6�P}P���~��7���ǹs��Q��ʔ��>å�fFfݔ�leՊ��^���JK���D+�D-�g�q�J
i�\�rT��?8z��Dh��(~BҠs�l���Ϣ��J$��3**�1l��+�a&9�$D�g���?�KY6|�T�՛�땰N]}S_Co���W37m�} �r㮌�ױ�1�̿+�F@O^�N�^a�:RV�q�!=i��R��nñߡ�"`	��e��<��&�2kn�|�OB���B�G�㞊�"�˚VYcQ(�_�Q��j��]gA⻫y���?B���f��ǧ�6���Q�&O,>�����!�TG =�>�����'5;�%�s�~@��P�H��o_����kg�	���25�Ƀ)����R�^�pd� ���{��Y[VN�G0��y�2	���|������1E�L���n��*���5��*yWm8u:�5��mV^dw �*IݾL����ꓡ,f�1vu�l�A�6��b	|��&����!�\%c��� ���?��+ ����Ǹ+ojA86�b�뺼��/l��Ob8�����¦{���o-A*�� ����8�%z:���6����/�|�M$���Qȶ^˨��D���7����^ǆ�:�3�+��*�Y%�{2L�~u�k�*⌤!^�R���q����F�	O�:"�w��Fɠ)��k�J}sٚ�N�i*�o�`�~�I��ݒ��:�Y�MZ:VU����7eH'P�:��|ӥ���1Q�t��JrX�7O�_�<�m���7 ����E�1M]�_�����ekH�[ڬ�'n��\�U�(f�;�F����#�R�Zzr����,n|��"LL!0��N�VU���u��h�f�;�5��.�s�g�eV㯗v_��BT�����92جM?�P�@E��8����Ͷl4!d��Ģ��<�y�Y~`�߱�2�[����K�-��$c��ݪ�ī%Zj{^����O�馢����ł���JX{��6��2_���C�3y�U[�t2ͪ%�gΗ7�IES{�Z^~A��
UF=�͋ĘE�bޝ��B���M��ñ�P.wH/�D�P�>"Y��Vĵ���>yU?����D��=fT�CK��u�:ə��
���회߆�/AK��D�~�g�j��������KL���yU��XD�jLU�0�Pv F��U� +�s��&�2|�c��j:��b.*2Uc�5ۂ�g�p�M�r����y�(��V7#WK왓����W^� ��n��H��_�����0�X��!^������V��sǜ���v��i����WV(��c�O��A_���~�]k��{����.�:-���� ��kn0��i�8aZΠ�&|�2�Lġ��S̷���2)��߁2��T>H���⫖��9�e�+�f�]���^&�I�#��yX;C½���n��OՌI��8׏���O=Z��c�γaᎿ��39G�,������矇f<���k�(�x�;x�]�vl`�dIk�TXH��e��}X���Z���t�M��X�ֱ����QL�U�Ӣ¡�Sܣy�}G�r<���.^%������T
Eַo˹�kl�V[S����{=���"*�|W�R�|U,�p��(J'�����r�z�N��S�z�p��F��t�۟���;����z��Ҫji�\_[@<�^�R�B)��@����������f:`�X��_�6Y� ȸN[�k�MJg����d4Ɨ�Y� e�c�.f���ԈCz&�����98��Z;�l^!m?L�h���8�
�'��-I�l��D�X�~��)�����9b�$<��=��:vDU*��X/Sda`��DQ��?2_>�Bүã��#5��.��W%&[���V��s���n�rs�7%��e3{(D�+��{�(p�'�TM�����`����sq:5�\������2O&����DGmf�e$�:���M��U�Ƃ���&f��5;�I�~��������2���4�1��6�*�"kk�ª4��C��vA:6i�3;�%
�ߛ�-Sc��D�o���܎�v��&��	�+x�V�hj���Z<�|�U.~7�
�T����^۶�f����,bMN�ۋ.y�eJ�� ��<��`\R�7����sҌ�ÿC�:;���������Lr�wC�+�����֒���s,��э���ϕ��l�Z���
��@�K��nr�P���sW���e]����E��Ӯ�zB	J�<�?�U�#�}Tf�x�2���h��[y�&w@(�%��ܞk�>�j$�:��[g=�"�;
��2�m�C���X7$��?t�4j����,����~�� hc���*�^)��m�G��0=�'�VC�=�����O�'���ap��ɤ�ⲭ�|�h��貏��b$���CC���n/�QD��%�ci8�*4��s=�W6�Ae�lIʷg5��͈vSr7+�۱�\+ft���?��E��x:�n�(�K��g��p��7)*L�e����+p��C�6���_(xైݼS�ҝ�娂�a������p�p8R�+$�Y��ǩ@'b�W}>��jW��o�"3l����/Z f]�)�Q�7�!�HR�֯I|b����q����)_"y`� C��W+VȻ(�2;{�$k����Z�3`�`m���4%�@X��|B�Z�� �޳s���{MD�k]�T>,vS�OU�ps˃��fPcHq�K�����;ޏ�jY�^��c�,��0J�	b`�V�:轴�/�E��<��)`������9��l\̮��`�	M�Z8ՙ�τ���t��ll��*� 
�p��<�X� �W���(��A�Q�q� O*�`Ȕ-wS��\1���;���-t�_,�{��ȱ�ҘZ|� �v\�,�~&@�/���0D�bz�D_(m�!�𱽸i��aw�"�R leo����Ff�K�}�&�z�����E��5�2� 53�sP���t}f�]�i��K������H}�-ȱ�L�]VA?�]�zB�,e��='co�g�R�s+��JP��HU����E�e��XN��,w���; �J�sr���^;�_�~�!�F���.
ϒ�r�^`Z�&+l���d�̩� �X��r��GY'��W�;�P��9�"�|� O�+F�4��oݢ���xr.M�s������Q�ܽοٳk"�,�EϾMT�	.���y���7�M��q�hl,# u3���Aђ(����7��K!0'{�#~�	B��l��o�����v�֢��P娖U�.�&��@�}�?�ioVƬ���_il�;F;���Y1ܡ�z�yJ^Ы�g���8��9�4]�� ;��R�a�E��rDGj'&���`}�$9��o�"��5�-є�v��y�� œ���mhmPEC�N�W{�rS<,co;�\�3b�hr$i�8~�˂ٛ���+j��M^K�od�ژ`B���i%�`���o�#�3��>�����.�e����a]K�1��*��f�)"\�� ���@q����%iL8�
����yg�{���g�7y����n�Z�A-���bo�S�ސ�4��b��
����Ʌ}N��� �<�Rʧ儍���O����08d�	�ub� ǯ4�"i�`.!�����9�(�����Ėk�-xk�6�M[�n�N��˿ ˧BhǝU�J��1�)��~������Z��GU�E��8%WG�PJ���[���\:���:���C.i#�({[��0/�\�!����S�UM޼ C*�!�<��J�[��d��$�X �"4{���yy�^����S`+�3�>�~k^q%�c��]�5�31Z�?�\q1���A���ǅ1^�iz�ό�fZ"Þ&��!:z�K��o=\�o�Z��R��r��H�֧���j��/{���K��9'	W��M2��9םawZ���B�Ƴd���l$``H�#�⁪��� G�4
6� %��l*�E3	���-�|��k��;r�cܳ\���#��[����'۲�W�Y�<�ޥa�Đ �eݿ"K+��s7��>��>suO	�g�K& �>2�Ժ��6�[��+�E�'��T�� Ww�Ο�c-o�.���0����gi*�ݺ��C�9Uѹ!�:���ě��/��(��ޒ+�&|u-��W��]����N�<���W�~M��kdo�7���"�i��Ԛ���-��\*�r/�α�ӽ;;D��[��V���:�Y*�@܃��xFuΧ�4��j'$95SaIEOVD���5~|�`0��rcBd� ����d��j��t�7�����	�K��\��F�[��]��{_Z��ɫ��-�X����^p����]P<��Una�W��p1^��ɀ�k�I�����}`4�+1y��]�yC���[S�7�Y���"�:?h�/�(b6��Db��ggөk��siK��HI�(Nis0ǜb*�5[(Fr��������I:��I�A���z����6�]F�@�I2+���jx�W���nU���J�`�9�?K� ���U��r۴�(��������|#%��d�J������FY�R2��b��վ�ſ�Jp;_昰�5�/��J1.wp<f2v�ؽM�ϐu�ZîLI����$�Xc��g������L�F��~>��W�MK�^΂�����Պ�SqW�z�O�i����&�D��Lk973�`'��R;V-<����(��R�݂o��#�s �R��!�f��~�09!� ����!���t:���i�꺞����`TA��!<.:�v�7�⌛�� ���j,����(7�3J��&�z�h�0&���Y�A��]���w��!̆͡
�'�RT���ZdW k���%/�=:��b��g%� ��ն��C�N�����p~�̄>,�Å��d�������a8#�]�L�LM�O}rs���+kl�缙6H�0 �X*��*B�i��:Pa�/�y���j�\3,D뫟]�$�����Lsd�E~A����hިeCY����M ��/ �<�Xg�d�
�Ig�|�>'�.��:�n��~��4�g����N� Die�Y��	c8���0	z�F-_%)=w��U�C��'�V(�	�y����K3NL���p��w�x��y��9��ä��ɡ�Lȱ���NW.;����:�i�n�xq��q���% �[�7QEZ���V��"�a����Q$�p((���D(<E�:�`a�A�0�� �5߳��h'�f�g�[I�S�Tr�Ł�qA�8қ�f�Xp
5���V��Y=}Hyux�_�p�#�?��}�vݍ!���"@�G�8-�ξ��ںE��P��0�j-چ���E�`�Z���2��=;��g*��\�#���~J:��'��=>P��ϟ|�b7����t���wg'̎���2��3-�/L�_��gI���̄U'�=�L��*}��V�C�)F�F�'�Ǜ�4w��2�E��
�����AqE[���aL`ɹ�tB��b��(I�z`�m9L��T�N$��M�9v�V��� �/Q�Sp��2�화�_Pw���ZӁ�Q2Djy`ٟ�W��h�.�VQ��$E$�;7�ǫ��1����7�t[�!���ŷe��:a�*�L����V@'`�вzBenf2� Q2�����P��t�Mr�Iff3������]-�S�lf�PU�gQ�dOS7逆��S.��1�~���՛�$x�([R}\WLE��~=f�\Ȅ����=a��VC˗]�a��xhzݚ�[�3PFyMKh��i�H�������+bY��?���
4�^�*�pO������!��AY��Xd��3�����$�j2i��@��L�L���̲|��ʰ�TY�x.�{z��I�H�y�4���&�
��Q񰽄z���&����3�6I"������v�m���'_v����G�P��}�0����9~'���p��I/gTjy��bN�5�/>�Qgi#5��5X+"���s��0���W�&�\G&)?j�o��,�r���AP���܊o�p�%��w���z�l�G��d哔��K���Q, EAq�Ug�o� �����v��{f�W.����@�[�f�ގi�������E�'�
������a���f�A���ԣ͢��Ǯ��	��X߇��C%
y�Oj�����@�k�lpY8�hS/�@x�ifѲŷ1/p��#e�,�X��?RQ�1��C�!��
��y;����dn���3��F�5,�BW����1K�b% ѥ�I��	��
Q��[w�П>�jQ G�Y,�a�l���w$����K��K�iW���'k꿋^��s���Qh]TG�MJ̤��¹�/fgL�	p�uWI��.��hQ��S��4����]b��v$Og�se�KA`TMfI�����徖�R �%j�dN�:��7 4�0:�אFN�}\Fj��Xh���
kQZܨ_F���.�9�de����˩��[�r�k�*(K�_����dv���P���m/2�B��+_���%5��a���®&L��������!3����b�
�7h�6����(����"㹙#��?@���HT:�sA��2L�R0��Rn5CY��)T�C��;���������/"+Φ4?��
�Bx�0jXn������SC(���5S� �֢djn&�L~�y09�_��M�8��$�
�>Y��AN�qW/#"dV�A�D^�����W }r!���8�������۱���~m�����m�R.��1��0#��`���u_�*$?�+�-�3���$vAi�JN�S��&���0���}�	/��h���8������?7I��4��ʾ�㪭뼫Y?*�=C�\V2=Ziή6h[f���8���Fl<fufm�U��T`�r���8ġ~�<0x��K�IT������	�֣�)#��0�^u������g�y�%���7�� >o���lA��̨ea��M�_� ���&�{�`�?I^ �L�h����L�/%����c���4��U�0�d����.x�����T�P?�L��`K'�}���eۗ��~��[mX�,�Ѕ|��)>M�	8���#�Y�sA��
�Lr��k�?�_h�ڏ��%���y�EiZ3����V��)20�SH�"��=�܏�袶B����h�]�t���cV��5b�� h������5J吶��bǥ!�c����S�s�N�����&}_�9��	�Y���Zkt/�>,߬�ū Bs�׌��:���;Z.����+]~�]�պ拡�T�)��1�2��]�ŏ;�M^����N�1Q�~��1�a�=�^8g�9�EYS��F��{M[���5���.f����<y�?���ڻ�8T�r�4ey}[�������AQ%����N\L���
�3uW+��k'��
e�� �"[ک�c�\�u
?�1z&���%]H��~i�?�Q�fK�� +jb& ��a ��Z�+I���2� ���k��9h�%^�@c�ʧ��f3l��?�8���lG�ppi��
��l"���pZX�1ڊ)ڝ�f��p��*�DW��+�+��zuC,z���Α�����RRK���1�l������p��3;��f�beZϓ�{���^��r���]Al�i����	�׭�~ҟ��{���^������l ����lw������9sd�i5u�����O}�7b�� ,���2)$��3��k������0�R��r0	nB��h|J��{=6��_�h	�4�K�&I�`�:�K��$֩�j���F�R����4�괗��,�,�)Qe��J���}��xh$�ȡ%�N�:hu
�V��ZMI�V��\����*$:d��]檾�m�v���1(��~_�ftuQKI��I/:�ԥ�Pܿ��f�1�y #����t������Bk�����\�r�a�b'��dqa���nf��L�$�Mjc�d��n6#�L��Ǒ}fw���b�\���01���<��k�奊98u ǖ]�������Gl&���n�ˋ�.X�9��Qc��X�*{}�6�m��.=�c��ޛ **A�� �_v�M&	����$ɮdz��?�?X�r�VY��P���T��9n�[˲i��tR�wf `�uR#sD˔�@�>;h>�X���w��=flL���|�[]QS���&�?��ɽ�VR��	>����*�#�e�L��m��92�I��v�s�7�TDL�R�ꈝAF�e	P�q J��ҏa.��V�������bFP��x�X��͝hcJ�55$s�UV�
Ճ��?Q���Zɗau�5�j��V.�J����UQ^�Ȳ:��c�W�]9����9�}z��jL=����������2�;�ZYO��L��4��Jz�8/q9��7��wd�ru}S�_ �c�W<���Dx`�̶Gk��vj��UP��n���Y�/�U��6�z�4w)/m��uщ�������$<�x��8�������{�ր��^w2�W��M0�T�K�1� �b�J<V�^����#N�eV��O+����DA0#[#�?O�}�0��W�|Ĩ�+i#R�PH �=Śz��¸�?��Q��Q���*��
�)�<�U�R���[,q�П|,B�����{��h��J�89�K">ݝ*VXZ��
�2�r���\~X�^��|��pX)���0ir�����0���Ǻ�@�4���[x�7\?�1q�RT����aJd˸|��,�a�tN�N9XnP�KPD��c���i�lV)���KB%�yIb��/�xs�sG�.�,�1��=!-��y:x-{�^�
z�ãs\�l���r<_�(�ZU,p�8�}���T�<Yt,ݪo~��1�?��o�hy�k&^�:� �
�Z���~0�-�LG��ne�%D���]��2q#Z_��U�r>�	�#���	�?p��}-5:�^o��*��6$���aˋ�K���Hċ����&������C�ާ(n���bƤ����X�>P�7T��>��"l�n������@	}gݠ5�p��l�h(�dp�㫏ԎT�Y}�+[#(��א�����T�̊��.��?6</
>lI.PŮ�Ęvj�U}��MIwٰjA	}������y�&�y�b�������Y]tav��n>E�I>�8bXv67�*��0�%��!�T��:Λ��'��p�J�ŏ'W�[���J�<�χD��-¦�Wҫr~=�`'�-��si���;G�_��X��n� �*팞�%p��[�ⵈ0�%<-:g�et&���E��'~%|�|�=���z|��� ����i�����[揁m;��Ŭ�s��J�ͼg�:lTug��۾��cH��(�Ձ�����D#wm��;+��{��'���`�~�����Bt��9��}�c�M�@�F2,SPZ9Z-�@�H,qҴ1��)�$��&ٌm�����jY��X��ՠ����@��%>��Q��wG:rl�����a�����秨��#O�����-�����'���jQ�*޺��",`�7{��N;�ͯX�ꡮ+�D>���*����z]K1Q��o{z�������w$��r����Ɏ[���g��a����Yv繁��'jk�)So8����@�#���t�#ej��#(��@�H����Bm�q<ȨI�o����,8�S���?s9�,u���$}Wj�̼�HfUB���'�-n ��?��r�֧x�O�}����Q���u�^'z�ᐣG����zJ��M,�<�#UP��,��d��_5`�~��N�L��H�w�g��Cռ��ۈ���~�z�N]��<���儒"��I�nFfH3�500�0c��8s�!�.���yYW8oF�9�7F0�"wܩ�����qԈ��,0&R0�	�ٓ�mj�J�����ҕ֑������抬V��[��y�z���1y�������*j��_��-�C�^��8�S��?g�3��n6�3�ڣ��|([g5�����O޳b�5���j�>i}��»��c�D�<}�9��!��bT.��c�������W��D�Og��Z?6�zKwR-�0�bn�ڣY���Gf�0Hm8����$ K�����C��O���Hh0����ó��?=�Wdٍ�XĂ,�&��~�����@�H�$��.1�h�Ɍ�G�nʳ�LE ����B2��?M�&)��-�x�;a� }���!�ʐ��n%�| ��m�2�`�-M)�	�/~��͡6��[ t�{w(�������5�7Z��LH�U��,J:�Ñu�_ij�iQj�hJ/��+`,~A�{��?J4��Ӹ�ZҐf7���[�)jG|�˓g4, ��HR�����1v�����B�
ͳ,-�K���jde���
ye<$N�l���Ё:/��
��[p��#DZ#�1n�+\��|��\��	��i��a�a]e&ן�#H���L5C<��c�j�<%���5�J�1��,_o��Eo*q�n�!]
���ig�m���x��U⊥cz�����F���b^Mb���aMP箶��.���y��K�YDbK�`Ar��B& Ƀn �f:��MVl���ވ
ɺ����C,�"������&�Vb|]�;�E�����t��\��}5�/�ڶO㲲CWJ��8���B\��#7� Yup�<�G�Q��6h����:Zt^[-�[�Dp�uYq�]�4�5��N�S7J��P&4�?�%�v���7�	�*q:�"~���O�O4O}�8��j��d,�u�������m)e,���YGE$J���z�JO{��|yZ��#0�5��X�A�2��i�֝搂B*^��%��.�
5�:���i�Z �R���-��L���Y^0�[̼\�E�Gi�����c0��n��%��:!�-	A��4��2��-���-��R�,����`伶h���x��U�Goƥ���55�ԣ8���p��
�vw�B�c����^�����D~T}�:.�P۹ 8U�
S�1R�R���u
l�C�^ڼK����k�i���Z�h�Hd.(�p��e�/�B�#����v3~m���?� F;��܎=�7���P����5�/��hZ�f���\gU��������}��1���͙u��	j(76ٱJJM[��Y1��w�t��B�#�S	1�Նa�W[����nK��=3������^��m�5wCC��UB�Xi~w�6m�搩��To��1Gh����"��oG�~n���t�%h��ō�8���E��a�{g�E��"Kj�.4Ơg���%��fW�4̑�rgm��ƾ.��8���L���t�LA�dT��#����*E�d��_E��Bꎖ�P�g�=�D����s�7��A�4�o$���8���w�.߅�p;��{�\
0k�4�}�j\0�p�x]P�}W�
���h���	����j���xo��z{�����u�u�H0br�jǯ�()�. �u*?�%���o��`yu>���Gp/�f�P�����D��O.2�`�J�I��y	ۂp�r�g�-���	x1$� �a��`����}s؈�AO�xlN�xd� ��Ӿ�V�6%�/��S0���g�Q�b7��T�	z�~��>��<���/e�����53`��W^I��
�&ؿ9�gЦ+�4��X�N<X�H6��F3��Y_��:L--Xe �ɗ{��S@��@��71���/��F���o4GO�"*�a3ŭ�PNؒ�	do�;��� �	��!�f�Q��7.Zڣ#�����������c�39�⟑t�c2�ά���t �-�ѨX��zr��u���q�#���x��a�E]>YS�\�5i��RR\w���ϊ=��QqToI?o�����7@��E3��2 �ݍ�L����ϗ[�,�_�>/ ���KRX���aD��� ��"\J�5ցv#�gv�x�i#�����K=�,�a8ƫkL�M%#g|��W�C}�7)�㵷��~�z��90hڦbΰ����~|9C��hʔ�c��j�"9GPUtp��#L[m��_�p��y/[<�	�}����X�e��P��C���ɜK�`6�h�H64���lV�9B�~�$�CU����sv���4���g~-)�׷�n��h����L�l� {��c�k��<��Iŗ6�F�]K�EkF؄V���W�1%�E �V�Iά�&�4��4�$ͫϏQ�P��X��/�'���b`G|rĕ���PSK�-q��	��P0�����@����l2���[mv�Q\)&� 1��s�#�"2u��|7�WW�����}��1k��L]�:/�ʙ�t���0��hptn�0����{�p������E�s�f�B˻OM�Q	���G���(-7�蛘O�
��ȫ��Ǟ�nd�x�U|n*�[�='%���{Τ�i>'7�sD2�h)u���.�E�}�"�s�&�&�*�y���q,�	��8�M�R�C{�GQ0��Kj�6b�Ú�'�$���Y:��J�m�ĥ����@�$�%�@*��xb{��-s.\���O��Un�_��_[7:�+x�X�����N��B���v:|��ޓ>�C��v .��B��i�������z�$BU���6���b�}f.�Y�<8B���F#	�K#����y�O����Qk�3	��:�]<N2E����.�1�����;�`>�7�Z�hDn5箨C��V{��4���<wc;<�T��"QR�Ox�J�ۥQB��q���:�8j@v���t� �����LH���nz\����w���_\�];�<1֤���v�I�h�����S<��5Ҥ]C|����_��vt�+U��A/����'�E��<@Y��`�t��]���5ׁ��|q��~$Î	���/R�sYc����~��ˇ^N��nf-�6���
*0��5o��3%d°V�����ݑ4b�FT� `�ٮ�[}��v�,���qiI� S�w�#�y]���:do���.���LD�w[�����h�PݿP���ǬFv��|��);<tV�Nٹ>�Ť,��������1|��y���E��ct9���lÆ&s�x�ŭ;���#��F,�ʋ��U�R���ѱ���M'/ҏ���v ۅ0��;�����Vrc-��!�>J�{\�Che����_�
(�V֍���4'���p3���Z�Ui,��p�;��.]>�� E�N���s�K�S ���iA��O-į��}��u+�E\@e)B.ln��V���Q�W�b��P����:3ex	�:5�9kR��������o���>�����i�E���g�@�$#Ҿnѥ��ɴ{���%�$�HGf[\s��0����\�3<r2LU���W��x��[��1 ������5;�p"�T��O���m�E��Hp>�6��9j˜��
��"�n�R�e,Sιkw�HȎm�̞��%�!�9d9F���M8ikޚ�x���xO�x�+f��r��zgn�4*��١%!�3�k�&��s��X����{�������b<�aj�zH�wA�輁�J[ֱY6�D=���O@��	�=����K㚗`����f��y8:�����Pg��#Z�1a��e��Js��B���b�槷"6cc[�[��^H��aXc�߁f�����[���{���~��ua|�+H5��#�p`�{PX<�� �������qg������s7��j}�0�	eڗ��C�������_<���Z�,@Q�`O�t8o�T�ɦ�X�{d�Fq��|@�+��ǵ.h�����\��[N���TQ�7�w�,��;Fd�y&��UcE���4�x������J�S�F)�[��}��p�oO�/ŝZ�&i�|�-��Ù�7|��e�x֣��׊8Y��=�� |e�o|+:K���C~��`�Ra���u��4eK�8ę�TT��B�py7s�==K?�	}��1����l�Xc����n?=�k$J[���B���>:�%|�'k�^_�;���
� x����ǋ�j�q6J��7���Ѧı��}��XA᣼L�OY��Xb0�m���9m|`�\&�,a��s�b��#p��sf�;��m|(l�p��R�RZ:?Ǫ�t�G�k�LԹO��Y�W�cs����#�Ƞ�S����]���9.��n�;/ri����x���č��a���s��z���V*�/1_�1v}{��Duk�(R��r��J�T푿�0B{��@�?�~'�q���Lj�h��A͝�^�b�v����{:,t__�b.��q�������I
�s�瀠c�3��7<��mkܯ�P5�~��$yS�nmӁ�jþ �Z���!<������>Gt}�)�eƜh
�K��iL�����*�O)�r��������d��?D�5S:!��9��392��	��'��Y0`8B���
~J�CG�5�P��yv�U�Ù��,�J^�����Vo�x��>O� _�X@�0����"W)hǑ�uAq��!�������D�$
cb�Pg3Z����-�.`T�[jE��X��zh_��ݒ^*J���*���(���Ɗ��~|TS���k?<��2� Lh~z%�|N��v@�*�w�'��G�S ��g��+�Pg&��I�^��s�&�:�k�{��[������0�N��|��[���Z�¯XP�\��F?I;D@4�U�אrvx��|;�<n'D!#b���,M]�ئ�����JѿL�o�'v�W�j"V�F1�Q"�[�#�3`��5��5)/�+�A'�W4s$���A���%\�J_����ip��Ė0�g�����4փs8��)���Hĺ̻��.��y��&���]�s�=W|Uyk���@���$��/���½Y��r��h�6�}�/9yqI6I��Ou�i����)�����V�ܬ��U��&�\��F���5W���y��r�>E0����J䚟��o��~G؍@ɰ�a"Qg�� �bJ������K���;v�O�'4JH3��PC�Pfq�|$��`�ѳZ�J��05�&4�-p��������㈴e�VhN#�ԒF�`���̝�Y��˞QPw��3�ae���2�8>9E�os��g&c��9����A��^@+7��4¸J��Qx�5��쥣+�Ѐ������^���Q��b�nc�{_&:��Ђ����du��6aydk�(~�������bI��!��F�F��{�')�c�n�n�6�a�ܽS���^��ɋD��K�6@��媅���n��jq�m&b�`a�Ґ�.ukǩ����s�=���Ǡ�6.9W�˳��Vz�5#R�T�b����X�r�����xz�no t��Q�z�-3����%��%V�e�`'K�kb���]z]Q.K �Gc>�\�.�lj�gYi����p��Z�	�%�S�� O?��%�] ����c�Y�l
�ɫ�N�X�$�Eo�F�N���G%��_ѷ�eh4:��t�`�XU��Q�G�� �N^�?�8cZ6:^0� SI6���]5�Ȁ:-*#��������T�.�$�6����
�=�|z�b�j�>O��L��H]��A��h&@��U�Y8�v�X!��A����`�K����$
� �xYa��]0Y�DQE�dj�E�����Q��7���I�I ��ju���Q�}�(�嫴H&qc1��0b�����=��2X�Bn2����h_3����C�0����>߄t�����*e#9���f֐�*�2iM�r�=	��n~)��m0+�y$��h�5R��o� 7���H��HNآ&)����M�.�@g^�lXP�^B������w�B������t[�C��:��u��� �_�w+	l���9���P�� �ns}fʾ�t��<���ęf%jk+\Y�"��o��A��MdX��$�����@֣�`��@�ؼUC�&Jh��$�-~<�s)4 ,�v{;2�ɞ�r�3P����u�6�>��p/R12��� �!Wtd�}P��<O��������Е@ &���I���Q^9�fNg m�a���:-�	�i���2��p�R��F�)�s�S�ٮ8G���{�cY��ڦ���-c7k`���w�M�@z���ǜ�:Ue�p�xy��p"��]a�֊ �K�vvt���\��	���O1o�%��E��!�>ț�����\�[Z2ش��e���J��q_%��$���R�u�`Ke(��sv�`�O�,�+�\Uw��t����'�a����E{vK�E�y2|~�_� TÁ�i�MH�ͷq�����F�ɏ8�q�9��u_:
*���05��R�Ǐ�����X�,?����-����#&��W?ϓC��k�����]5CI$4}�B����pz��l�h�j��0�]kD��������0�)�[|t�=���M�<o8�iݔ�X��)k���ֳ�+�� "���kU���<���pb���b�����������"�s�..�N����6�:�Oz���
@zY7��ZTCP��@Rs ����R\y�j`V �] sN6d@����_p�ͷvj�+��+�T�#��pBF�¥��NjK�ª�睆�v�^y` ����-58�d��4	
7X"(q$Q�6z�ȶq6��g{ �����fM�Ed�z�φ���6��(�x���3�8k�?T�_d�o�p/�9\���z�H�A�/̽	5�o$ �J�7�gn���w����|�p�5�"Y���&��x��1!�z@�ĄC�� 61�;K�K�|b
ܷM������5�2X����bڕ�]2R��e'�p��Yu���g�i^�����;��hjmJDo�蜦����i/B�0��b��0�P[V�4$�nX˵?������m�]5��Bf~ի -/I �t�i�w�-Zz�=���Bh�YB��_z�#���֎��6'4ɏv(�Ua���j�+��%;ͣ�ՙ`2��Ō�xO��'��� }ܡ16�ވF��ʹ�p
�q��<��S���3�81�p�:�,��w��{ �sr?f���$�3�@����s�8	�b��W�n��b
��Ԡ���</���v��*���5��\�d�u(�|�N�7h�&z�5�M[R���V{�t<�ҿd\����L�m�����V�]\�Jʩ�?���gYܗ*�i���w���/7Z�2�p�����t�#�+��߉����T�x.@�M1)�O�>����@��Iؒ��otSYO;nCU�����LN���~�}�u���.�D�}H��ل�>Be���$9t�ל *<�w���ѫ^�O���N�0G�<R��D��ٌ�^8h3���9wDSw̞3f��L��ѐZ������nW�\(Db:�g������m�HϪG/�Dm��[ʺ}8@�ѕZ^�^��e��{�ix�W�y�u��#~���do���ÁR-zx��F��A��� �7!q79���IdQqU�� �S�4s��q��89:�L���	y�#�^/�~c6���W��p%�j_�r�L{A�
 <��*���_d	 Pe5���c�!'��T7@�:u�S�Aq@��P�������Y[d-�C����+o�[��R����C�4����O~��m~��J>��{l��)^�%��1��e<
���f	��sxE����IetF���=F#%��牘�b�M��-�v$�ہQ�b6"��ɡb�yv��A�-��"3T^�+A[L<�|ȄùΑ?���Q���b�W�%� ��<��l�t����vi��kD� [K`���M���l���2�u��-t����˪��~NbLڮ���$�"�c��a����r�Y�%-{�~��@�\�o�ǝ�oG#��Us�;<�B�ܸc[*��n.:�x�o����j��1s>���p��n�?��Ү�ZHe�44��a7�9я�0���^e��wv[27%�C���u>��^�-\�S����ɯ-��O
�+�G���";!�(�2?���#Zұ)BL_��|JP���WΰH�]�&M��Q�s�}�/�Puן'��0�J��N�Igh�^��}�1�;�\�S�6�{�r��������VjI�>g�׾�DѤ�kk��do�3`��PɉxLB:2e����^3+�3�jV�乐"%��G���p�����B��)-�����9��1<�S��|`�o�ߙ{��n�QE݃Wn��)��0p1jp�����ì��y즗���3y|�F�V�q�������R����%�#��>��p���p)�zB����A�hLo�Ǖ%B޲A���3 |���h�Kbb��Ӭ�Bi�`�?w$oUY#����J�:�~�yp��Wm�j,�O�^���tt�3��T<�Ҏ�C�,�a���1ôƺ�򳡽�B�H�C��n��	��6��)(�!Z!6cN�Ɇ-W`�H�������g�ݪ�h�W(�YsT8�c9U������nN�;���NU*˂�k�
�'��B�����D�e���~�k߈�AnU��6����~���BCM�oK�d֟+����U�n#K[Zg-�إԧ��F㳰2��o2�4�.<ȗ���Bަ����qr�p�5L���CH7�1?W��}Y&�-�5�P�J�e=�/Y�7�O��-���4� ?��e�b`g�	(;{���ZT,���P�&)�@6��ۛ�9JJa2N�'�,�:n�i.4W|w�M,q�`�%�.�O� � J�Io�3INP�1}��
�b�>�����n����<���<���c��!�I&������VNx�����ҭ�2x��rW�k�.�!�U#�����\SLzVic6;���]A[�I�'��`�\;���Z8,�T��'�vʨ�p�#���ۚ<�׸)җ}����9�����Q�����v�ŭ�s�Oʵ��oG))>yLv�9�>Zd��S�~5�b��x��B�j�O3_2�9g���ȟFS�H��U�%V*�@��pdG�DU0�L�;X����콌#�)�czH�]��T��C�c��7����A�=$�~����q���fp�����1J6��h�o�RCc�����G�Y��^'Ɩ���7�u��3�C�����l��㖹��=�g�/.��������$�ԓIj����b	Q��L��Hz˘,��)�9�QE�����"[G9��հ2$JE=��B�cE�������by�"�����r�����<�oĜ≉>��}�U�9���&�.�ETB	m�_?��k'��[�w�h%�#��˖�����4��M�Du��K�r+���
�	\@�ӹ��	[��
��n\WLcP>(כ������G�u6S��E�������@�[	d�qrY�X0��k�G�T�����7]Awr��n���d�]B��](y�~�ϫ"M�c�yb����\�l�x�8Q!�,2m�C��f���&H�e��z��I^M���`��R�H�U�1T�D]����6E
�3c�
TD�2�?+O�6�
R����,à _�ޣ��8jh@�Yiua����e��Fg.� C����^�HV�'�h�ֵH�=���^bA�B4A�?yrMt��"����z��3p\�_U�!�^T�ؔ�K$^dC)
��ٶ��ge�
k�+�r����	{�]n��T�F�:Y�������C�~��,�-1b��JlF�lM����2Y�����+�Dc�œN�3j�}�8��7����=��`�]����靷+f��=D3������歰Oo!ƹ爝H��b�
p-�p<:�J���P�~�:Vrz�d?Jtn
QhU����#�3*�������Ū,.��^:�������gr��LL�,RUHtb�*j|#0խ ")������[d�E������;��ۣ[^�0k\U�]^d�'ǧ..S�u�$葯�>���E��w��`L*8�.�g�q�zb�9#�%#1	~�E]Q�*�i����J�J��n�Z�����F����{�o��w�D�>n�B�L/�D ��g����SU��}x�8�� t[~��P��r�żl�e�n\�|�fq��b�^�@8���1&���;��s��p�����¼@_r�Џ9�Z�������D�7<J�����R��p��+ڽ9W�[��z�1�b)ж��/JM���
�Fڼ7���2�<}#���[�����ޣ~�_{oQ6JQ�ű{b
�� B?s�9-�S�>�����g.�c�7� ��_~Ϯʺd"�Y�ȱ����AJА�g1������Y�p�R|"&TѕGs'�Nc��Fyb&�\d��Q�E �*�x��<Ε����^��W�Z��#h�9�636�C+�g�L�Z��Q��?�/6�Y�'T�i@�١����OȮ���8�N�N��|��|l��/@�}"5O?yb{��1#��L#N����s� 1�r�z�1
��V�C��X����&T���G.�f��3rD�A�Rƫ��T );%Q�K'�k�/��Mt��}��)E6���]�)S�,�ۂ��Y�g�^���f����pd�!hF\:����r�&�o���φ�BAg�J�sJD�n�wp����\������b	kZ/��6��_�M����E�/�Ҋ����Lߵ�b0��eY��EF�⿈���\��m��7q�*#�~����|��#y�����)����?k��m�W����YhL�m�vՂ�TL�ޔ>F'����d��0:���Qʽh5���?�ђ�����	K���m�JY�hS� �����\||V��tj�i6g
m�N���6�oIr��������Ξ��3�Q�s̐(��@J�}4���F� E�!@v����x&���7��C���5H����7�����e�x�Bu����#����3�l�"!�s�U�E��}0�b��P�\3��޻��k)�/�� ��j`R�j >-`g>���27}o6�^X-
/ qUb���������z+5�0����%N�)�H>�j�U�BD�E�3\w-��pi%�����h�W^}>7R�/�"p)`���4�SUZN}�lA5	�K1��^n���mgW��+seuwV
�,�T@�q��<��3��,8���rچk�F1�d�*�8���T��0Z$4�	6nBJ�,S�2=Q��v�~/[��1��;�{Tar*}ǜ=��n�V�ޞ���3|�:QCϙ��
����6�g���k���������|��\>�J��g�h(�U�3�3�0���:a�Asf����.��Q+K���k�M�J���)��3�S���3�vN;�l�xgM����Z��P�*��Sf�{$Eu�g���v�q���bӳ��A!?�F��D�9�g[b ��.J�����Ɇ_�t�%�}���򪗏&c"�m��^��* �����9mp�٢)@�b���|��_����f�:�OG-@,B4�(�����ؘU��ɢ>0��;��Uu����`�^��$��$�g9Gj�%�D��(�z��$�����f-�],,L�_ڌ��a��1<�
�Φ1�:^��m�����a���ټdO����FN7�gut�$�ؔj'�/�I�m)�_�;]���}_�H;����b�:��l-n��H�!Z?���N�K���L��Ҹ1�k�p�U"//0�c�\c��i���V�p��/�a�΋`�V7S�i��.n�4��aZ7�$ڞ����籱�6�$�C���mQ�Ȝ�c�M~���ԴP��/[��(�#ۇH��>e�܊��xֈ�[���ԟ�i���n1�8,�[:3"�],/]Ӝ'��=i�B{q�ab�x�Ɩ�鿼���[�KЅ�gmS�Ob�|W��)d��ײ�i�*�|�|=&�N@x�$K����:��|=褐U9
\�=��ϥ1�ZM�|��SҭA�e��d��nb^�U�ռ��>�5��`�_�ﮁ��~& ^�iCU!Vӆ�@f�I��>������֔��
����
@;���U���>2	�!ç�:�Be'��@�^0�nʭ�\��r��z\�S�9���;;�>l��{@�^?�j���� �w�)*p�OdS'����j�|^�Pa��"�0!F
T�qP�k���L��AM�R|��Ցx6�̠d�T�;u��"�q�0�:ِ@`���<��'z>ۡe�9���d��f��V`�����/8�O���.rY��»��L��l�n�2k��_qYdR]�S�!jj`�M� �:�nP~�BZ�����n^|1~��^V�ٯ~uK{W�*�y�-��ׅ�ԟ?�ק��|h~�vʥ�����Z/��ʉ ��
@CL	�em�����c��������H���Vf��+!������C����]����!U��v�[$!Eū-�Q�~u��D����{8�Rb�ܐL�l��8T�Ջ�Tƌڭ6j
�}v��?� ���(��,˹��s�N� �L6D�s4��C�����F���J�.�GXE�'ա���qi���%���}�\�w�J��H�����Xw� ��ӗ�4�l�3�{���ܸ3��NQ���K^p.~�9���/M��(G���2���=RS��ɭ����.�D���ˠ�)�s�_c�@��\�[�
���o0�G����X]D��	ZY�}ȷ���^�vOF�br�/(#Fc'������;����6%��߶���+��j��M_�~)Bj�'Pd��SRGT3|Wm������Q2C�3�d����Uz�Z��fľ᎜?N/�>*���=.'@��kem�.����D��s���Naw�WcӪ�P��Ntg��:T2-c�#d���O/!� �S�^��mɬE��fO��$~[ǌ��|-R���z]YE�� �5�
C��h�;q��W���!`4Wh��r��2��K!I����E����.Y{��se؃��B�T�n��zvPD�b�/�WM�jb�C�Y#�,�<@o�T,[?/���"f�Q��oZu[�9ǰc��al�x��K��ۄ�Vaׁ?��&ē�ډ��iKS���=ˈ���� j�\ �	�����(c�1g�{�%w���
�x���Fi��Ú,v�3,�>E�Ww���]�6��-Țr�)�$��Y �)��<O���SbN5�!툆�R�9��cj��X�M����v�ǎc4{k $�#�Y�e��(>�K�B�I��I���N�u���Rp������N��eԌg��F�5��]1��qŊ@o�F(�H���_]5����A�mK���ae���y�A�뎚kk����ew�\
�0 �p�>kɾ��`^��Ǚ�?������v�[1��yfQ0-e G�B~Wu��&�zE;���mf"#?��umK��`}G�fwy4��6;��v�(��P��dX��S	���!��I��;)2��`o��<��9/-q�F����}�	�Ɵ�Lq�P���6��\��dw�����l!MS�н|�75	Y2����m��3�P�%1�z΁L��R�AǑ���=|�����:"���o-��t��&�^��O�LF:xp�M�`=e̋Ks&͆ػ������f��m�! ��4���V�@�Y�(6��e�*��HV���ۅ#].%�P�#���;C؃�-��KWa-��Ei��sβ�!�-��N�'*zI",F��K��j��D��e��6�X����΄�,�:@L�׋�4=�F|FLjK9�n�����K�o�T�����uC
����X�����n���9������<LVC4a�}���,�mr��8c��i@a��a4h�ME�n�\o�R�;�7���nD�����;f�۲q�	o��`��B3��qKN7��-��Wԇn<s��*컼�1�M�i�}�8�'�/=��Hn��hB���?�Z �*^��'�s"q�JUnp���"��8�6EM������u�g�~>8�l�K�����E��D[มT�ιelL*1c.	�,�����<6�j�\oY�z��T�2��>�-�hSE�/����3�g�V;S�7���Q�'-�0��U(�ou�r�^�(MD{���n`)o���HK�:�z�7��?�}#a/��6�E-��/$A��R9�&��[ц�4|uH�:9��5\
&�dTF� �5���������ͻ"Nw�m��2~%��{�C,�_�����B���� }��$F	Tυ6���
7�.�n
6��H�R>���*y�7��f��~x��$�����b�3��+:X7�|W*A5S\Ѹ��L�᷶��H2�u�x=�V‣_�3s4J{TT�X�h\�������z<C	I�@R{3���|��^�z��/�d`�b��g�Yh� �u�?�q��k-D᲎����ř��3���rs1�w�O�?[��mM��w P��-�:��LT�[��҂@���Wb�t������3��0b����Md3�?Р,��7C6龨���h���/@�ej3⚪��6�Ou�,��m��4�	8�\� �o�����KvJ{j��N��X�)��E�\���CI~����2v��+�:H�H�(
	���aH�Pj _|�#[�Akr�m�5B����l���h|�Hs]�C��2���~K��_�	R$̘�3SsD���>����9 ����&E������A�]�!p�[��v&h�u�q!���x�]e�G3�|�fĝ{o>|���RI����[��<]��S�\�S/{�-*	�_���>�OGZ�_u��8gߺ���pn5n�ɱ��G�4?qMI�(����vi�m�����ج�-�p� "^�C��#�u,��I�MUeu����1$I�Va�hU��>k��A�f+�a�����L'�Z�F�i=��w�2a`�K�1��;6Ӭ��e������f3
P�$�X��q>n��2�͟��|����T��H:�C��)��)ý���VF�����7����<6�_8�2�a��S>,�'��U�R��Cd���Ȇ��s8���Ƿ�2�w:�-�l�#�F�G��>b���S�Q+�{��zg�U+& ����P?�έ{�P�q�~a���ޏÚps ~�/��g���E9�Ь��V�>���IUi;����:+p�=p��p�J��]��;/ *�c�e��Agf �)O+E=WO#Qj�KX�Ȯq�F�$S�.ɀ�&�r��W�M�I�fR��<A{�JD��}����MbQ�!�oxw�7
#�y�TH �6ή�� i�e�t�n�y�z�ɲ�*�3 �H���#��I�ڬ���o���
���l=�gBwU�`hb��w����D����(��&��ǫ�<������8m���)�̞U��s#�G:ʶ"T��� Ֆ�5f���Ó;�R��SԢ�S����Hư�$q�)-�5p�����mcq�vWчz�(]�[�f)���=ѸK���LL���y����Ъ�b�Q�=��	i1��2�C��3<��s1T����i]�;26�Ӓ!	ً�b~�V��TU}L4���1�%n{�!C�f��������v�\�[Z�O5	ȻM&oGhL�b"�-��΂�NV�hs�>�*?�ja��G;]��n���h	#�����Y��B(�O�.�Iʸ�
'X-o.޸�%�-�����6��s����n��)�Y�^i�;��t�X�B����(�#:�����tq��YTcҐ��/�&���:Sn|��/g��1+�8!����L� ��s������I\u�����뛫f�Y4HC�M���$����H�%�B�2����0�H��h�����uH>���k.�ګ��k)ڶ�z5u�01+�KZ�Q�T(��t��ت���g������N�J����Z�a�kv���5=�UD�X�*��[��:��1a�%���B䶛�N��(�x��ѡ��9D@2�(9AC����������d�ue���� c1�k�J\������<S�'+&���4��h�����'|ࡴ��X��\�_�@Q���Я�����6	�u��Q3\Z��5�/&=��^�x&�ǪX���Jar�/���f����������!��H�WKM�6�%?�;
Y�WRo��l[����CT�dp��6�0���4�C�渥{/��u�2��Kk?2ךw���|�S����*�v�j�!��%�s��h���Y,�D�=�S͘��
)?������2�s��0F�20��IU$ ��^�O<=�����*]�yoQ�gL&{=TNɤtH�w�ߖ�֜|�>��\�5!�z���A[�>��=�a� tTh��j�vu|8:��7��[�"��]���T��3�b�A�T�b"B3��N�lmT6�%T����'��ڻ	H�ł��=�̀ër�6��xU��R�.�؃ �O�>�T��t6��YP����N3=CT��ə���7��lMAx`�ڎ�;���Gc�����8y��Cm��8qcP0DF�1o����	��"b�8��Tr�{�1�C`u���Q���-��kd�����TR�Z�q�����6�	y8�xh�l�����>�8������<�D�Q|�6�ʟ��B�E�1X�M#av�ǰۧE)��0㩻���h������aQ��𔞳��
F�\�[�G2�G$� ������4�c+�[��Qoǁ�<��ɿ�	�`���pعÌ��ؼ±P���$	1��M���V����5� $�ZT �[ �|i�Д���}����А�r���1R�D,��:N��->��lAVI1ZL�'����xg�W� ba�(a��UϽ�����o<�2��� ��	6�j���g��í�Z2���(�{�d�.���`M����U+�_*<�RA�?��F&��}���]��� ���үy�Zq��N)�s�$��4+�8��bE�x���94?�IA�j��t[�\�SM��j�[�w%�`�E��'�
���HP'�ubA�ޓ��j�I2[)�b"I����pv�$��������gu�;x/~$�P�t&��f�Pļ���¯xt���ru��g-6��}�����'�8j��J4�Kn[���Z�D�����'ht����#��z�����Y�b�Yբ!��Ե�*\82���=8�+�R\�$�{;m.v����f&F��$�o�N�m�GqAL�[�Oz�:������ިZBGm������H�}�;q,Q���s II
C:T�AF��/�����W��Vs�"t��y73��m ��tqT�'�ԟt�2d�ß;���a��j��.??,�h���.0��y�i��~u)r`UK��dyh�Y�{�%A���Aԉ~���ᬜ.�O��d�/��H��IZ$^ez�x�j>�/RJ��<y�{�|������г6,���.��&��	=����f�njCw���yAv���UQ�����Z�Z������&�4��R�3ns�>hr�-+�&���+�f�)�(�+��ז��12��	!������C>��v�cvgj���1s����(�h��@�� ���Y�B��HO����tu���	W��K&H3I�I�T��;׳H��l�/Z�/���޾��۩�2�Z��b����77 fPC"�K�ŝ��=������?pbn8v�J�^t�ܒ�����H����Y)����'%�/
���^�m�� )S�/v� �J�0p��"f���G:�Ð74N��%!`�KX��]��tܝd4B;^F��!��(C���������t6��/�\?�eYD��"���<���j<?�;�/�;޻}�D�n�B��[L21�tBɚy��i����(r��o7|;�� �+'����u�fF�}��G��&Օ��u�u۝�^��Q��Ok�2��/�Gr̸A�i�(�@�>���y4Q��6�Ym}\X%]�4��R�gπڻ��y�����D�+d�R��\K��*U�w��J��y��V,Lv���{���R����1�r����Cĭ���C=kL��톫�:��Al*f�,h/ʕ/�F>o,N?��]O�T�U����[���Q*��GK�V����Q�����e�/b��LH���|*3�}�6�	��@q����!���$�$Z����a�)%���c_r�(��5�͏���).ս�Ȼ�+vm�u���E�΂"����M�_\,���b5Pl�<��NC�.�*c������v�Cg��2�ȡ	���e�LW��ʯ�!���1���N~��.�*�`u.=���ۥ���7�OX�é�A#�xi �̘:m����6s�|�>���ڱ�N��������pp�Y�����i@��9��l.F8\����R����6�V:ݘY����N:�I�.�p�ke��LW��S@��	K��1���V3	��\����V�NN���6Ѱ�y�=�\�#;X.1��'"���g:O�s�nU���5HP ��M}�:#��E}M
�K��AG^Y�H���R��F�{:$_ (��9�n�8.d��F�V.M99gD����[ތu��1�b�/
��$�c��0$��2t)S4L^J���<U��|����tjG��qA��>>��tI�6�Y�%�!e1Xd��P���^̩�,x��w
��R8��7T0� �^�iIN۾�NX ��&G7�R�9��be /#Y��A�w�n�#�*s�R�1G}j����|έ�q�^Թ�[kG`�*�x3k��Krt�&LY���%c":Y5���i��֨o�"oy��4�En����%K��l�&��k�������ۼ��1%Hdb�8}E @����T�#�h	���)��a����UG�hT�+2�(����ْq���!�ˇϐP2ȳ+}�.�4b+F^�`�z�%�V��u�a0�\-���e����I;�LA�(TrP�(���#=;��� Y2�� )���ſ���\�S�����KF5�gI=�'���<�J��Q#}D�H��A���ȰC���	�ȵ���H���(�h�߈e^�K��`:pW�i���2S�9y,#$Z54r��!wNE<��A�d?����$E����1#m!�V2�P�Y ���5�-bA{��	��ǦCy�.;�:||��#�[��G[/�;ާ H;2���E�K��Ǥ�]G����H���'�qa��0G:��1��)�p�HyI��70{]g�8�P�=��>�%R��a�,Q/=q7:�߷���|Uk7��PP}#\����χt]���?�ZY0���(Iܣ�(�=�y���d��r�R��b�Y��C�+�O[�$�u�����K�G��ۚ�Ϻ�҆��������#׼���i+1�7˚1(��I�#�Ǩc��G�J1u��v1 ��P킩�Hp�~���ٱp8��T�_��)���4��V�Ö�Ͼ�:�:p��&�%@��J)%���|�a��hX�����'�@�3&����<�vQ�&��CH�c�P�SC��E�x{>A��N�Z;ᄀ3���K��6�����;`U�>��gz�;�����|�g�)���t)��c�J������8>��6��=A__��v5Z;���bRӉ�#���BS72�p6T���t���q�f��[L�Ϋ�BlA�^�D��]�g��n�$�t����� �n���K��>��<�iC~4� ��wXH��f;���)3���uP��!F��X�!����f�Y���`������
/W�-�h��Q���D"�2i�w]~Ѕn	����HY*�L��N�7gg|fc��o�*Ud�ǉ���|�o�o�=BN�1+!C����D��k�����WuL��v���NVCM؟kD�L��}y��+�Ɲ&֭"���x3'�4�?�}*���/K�n�y���a^)�Sqsd�O�(��u�Yoֽ�ߧZ�4���{<��CK�t�����9���=�c�Bb\`��4��xq�58� Ka��b��(��.P�	M�oVW�4��P�;;t�Z��2�ea�&[�ZU�S��5�R��?�oÅ}�Ճ,�s�;��`�
�P�K6�k�͓��O���=uֶ�$e���p	P��B�;������3�:Z���|�>~s�S*��3����`k�\F�Y�q�m$�َ���1 ���E���IYw#0#Q"O
��>�u�	:�N�2Y8���<b�fm�ca��48�?�S)���_�3t�*�]�0�H�-F�z�h�pRؠ�%����8�1ۈ�~���h�5v����9�N/4!]����~,�J�zW�.l��z)s�mj�͜o���浴�7 8�<9�<����)������4Ʊsg��0w �Y�+����d��)�,6&߆�$�l�����{���K����WG��Lj��t���S�-g�: ��B!6�Ŵ"34�㫘� a�ЭζZ���[K� ��R%���h���]?��3�a�0O �Y>��Fa/�q�M���=�n�\Z��_V}��1	�Sq�5�2.-A��/N%��"T	;V�l~��=<��|����a�)���kH�)*������ / �,`R���|�Mbu����841�<�g�J���i4�X��:$ x4�� ���HQ���c�1���߻����q�'������J4��$,�+�nY�,BɆV����.+3�oJ�ӛW�^����@#^��X��Y��
�P�+}u%���T#��ܾ��ה|Cc�9������PsMFL6ỾY�׋�n]q!��f�"_�W�G������U�vj�O�4+:Sxe~M�p�qU�*�
���\�x`��R��P��$��I�|u�� �J�L�n��QxJOP�0GA� M��s��e���H$�AaŠ]8\O����:ߠ�Gl�U[]�b,��ix�hp��#ӱ3�x)�<��$M�f0���CR�$�d�Vi7ˠ���v�=,�@�B�񒨔��l��l]�N8!�j!d�:]�V�ҩf�i��l�)�>�J㻥�l*��Q4�jb�t��Q�eg�̎_�:�,�zQ�J X�5���#C��Gw�a9`� ��o�i9ypw����޶Cda�
��a���|��&
$���)�]����ĵN�-EQ{��.N�j��^X�Å���S���r3����	��h�0B<�A�T���68��t���S࣓AY=	%��"��,Fo�t�mM�<�)z(��1��փ�=}V�!�"»»�ET��<�tI�HUI��%4�j��ɢ��L���_���S0Lf�
�B+u���I2zDi��'ë9��ʆM����|H� ��o�^���l���0��px��)1�ҭq荼Z,\�ˇuZ����xY�EY����l��*3��(\!�����ֺ���=V=h>{����_\E����d��]m�Gqr�,�*��j�LX�t/���++����X0xU;GhVJ�W�)���w�[�]�@QR7O�+�p���F�a����������Uo����9=a��
�ت�o�����:�����C7����Y��c�T|_
�n�Ó=ó��� �௓�f"��P�}u�MC��4�
τ�H��D[�Фf��/��4���$�#�8��5��c�a�9��ٳG'ױL.RW�.Bm��!EsZ#��o��"����x�H4�)���'��Pi��́7f�1�Q��2��d_�Y��r�`���ָg�`3=2��H%gʿдXM��Y�[���B�r.�T��`S��vma�7dqD?U=�4�y�C�(xψ��mJ×�X���)�z�Hg28[��L�6֛:�T�A1�bm��Έ>A�ͻd2<ʱǫC�v)�����jc�S�`�=|�h�w�Dng�R�?�m����:bm~�&)ISap���r��'�բ2���N� r��^��XԊWϭ�x�#�wi��:���7q�	�ט���0���OS-x^�s"� �6�0���"<�G�� �i.��H+���]����mn�bo��%�P'ȼ�=A�s�-yQ�#�����y����5�Pi#1��G�)�'z!?�M&�Q�t#&���{w}q�S�UmHoXRH|�6��p�wl!�B&��R�Ğ����5����C��]@,�z����k�f� ��xa�U{��ukȉS�S�?�,'[�L'��H�O�}p1ܦ�'mΦ�n�m�p?�?JS�N�IK��:�!M�m8�ao�D	�g�9)=��Q�m:v��m�}��$���lk��XQs`����OO�ax`q��ZXV�=2�gq����Y5��f ��d% �W1lK���úi�`7�w[�*�*���r��Ul�����z���!~;���J��dC�HR�?w��(i�Kim�L�-VGzyY#C���$j�b��̑1�CϞ�@�`���Ҳ�M�%���-�bt_I�FGv�-�}M-���~��\�+2�]�j�Z���1 �UF�U2��UdvY�b��ޥ��_ʂ�MO}6g��TӺ�lʲa"�\������Y���8D��녤s�iDa��}� *z�UH�m�-�7�{�{�������Pg�c�Գ����<mO�S<�*FnG6�d�q֎Ѡ�|��0��tTr��uQ���]�^AgHw~ֺ8��Á�_(
��1�d�5��s}��cCEEπ�I���ӡ��T�H��F`
c��N�	0���d�uB��	ۂ�ܰx,暲{6^�F#�@��h��E����+�,�/�� ���\��}5���`~y�9z/X�ִ���3��2���]�����dO�[��<�-�����;������#��R��� b�t��ёE�H�i~����*�)k�s|��bw�6t�z�܌��da2�����7�{�U����T�~��sb����"�:I�׽w����ѓԸ]~�?|s�N��"S�'V��h��ܬa7�M��d�Vqۻ��|f��z�y��܌ks��a�jH`򕚽�B�JC���"�`��#5�8Žǌ`�:���T�x��Ϸ��g;+:��W0�Z��@�k�����0�g�/`N�<���� �/I��/�\@�V��Ld����! J2���U��ԃ�l:�1�r?�qU����|��R�$����|��U�@���ȹ�}JBa\����bo��C�hfx�L�q܆���t�kڀA��EF!t�M�I9oD+z��:����ZX\g��D�0h�F�����:�[Tt1�*��uԋ���#�r,�����]�q��5ë;�4��v�7AV���~��3�Ԅ���D�ށ�TKOG��Y?,D��NOJcZnv�H�_w�(^n��Q߹�����f���)͵֏]^&4z�q�9f���d����BvT���w. �i�v�0�����;q�_+IIg޼������z��>phYÖ��}(	�s�����v|}�� �T$�wZ_v���b5�n5�ɚ�j�ms5�{�X2�-��u/E^Q�$$�]H��Y/�. �V��Ȏ;�$<�w-��s��F���i O����k0gGn�I���OF��]���4I�y���G��C���v�C�\�
���:��)EL�/Rp���ab�Rh��m���W�c5+�ag�Ŷ2=�&�;;������cR���l �5���A��qV�0A���nE6�:�`Յ1�kCr��ٴUt��p�Ę���%��\��g���W'��eA��ϖk0��$䥁��.v�31o��D�T�G�Ϗs9�\��pzpO/�ߛb��'���۴�
�6�\WV�_p����'d����s���AFd�,�.�{PA��j�={�	OАMԬ-&�H�V���є�1����!TG���2���֨E��.a�	k�)��D?�MT���O�+�ó�l�J���g�?��QɁ��.T[�W7�:�{��Ǹ>��X����7u����א:��SGn�d����F�Ιr5?�ZG�'�t�@���������xWb�r$&��c�>�`K87¶6�~R���k*4���eo������K̃S���I�YQ��vC�m.�1��� Z���7`d
Apl�R/�̈�%�HQ�὾�rOͦ�X�v�O��˞s!þm�[)*����8w�8��VU�v����?wԳj�o���!�.s�%��D	Ad���|���6��0����o{;��Pf+�x�d�MEN-�����7�tT�U����ܽ��F �<B�C����й%iE69���s1�j	o$�A����Sq�Q���a�f�*���@������eB-�Z�f�"�X�I�v��{V�1o��yW8�Z~o��.�7��>6�vߊ(o�˗�����G�axw��J}�Lֽ�&7�*ڗ.�li��Dp���w�W�*:�嵏�@��:��_S�t�D���B�ЏC��aj���8
��'<,�a���F�X�ؒ���o~��u2y\�G�~�d��F���?��ӹ�CȡW�|��M�%��n���Tw1(�t�gZ댷��r���m�-����+	��p�Gو��(���if��4B��3� mD}���q�t `W��\�}����ڴ�[u��z,���H �v�4��Y�1C���#C�S���?� ��ṣ6!t���^f\5B�U��~��5��<7xyj�~�Sg�Фr�4�t�y���c�;�⒭��%�.Gɀ�M�>&/|U�e[���8�-Ħ�� �	�����%�Ⱦ�oR��
{��Զ���N̝�����I��@��x+��4̪��;��/d�%�]R��8����o�}|\vJ����Xn7���<\��oFm!>�s�.�8I���j�����PWCǒ�(lA���j�U���P�ɓO�^8j^���qd~�k9M����s�cJt��`��0;��b
%��E+{c!�=Ù�C�چ*/�<V�$�֫��~3�H�r��޹����_E(�,�4IB�f�d5���Ԇe��e���޴�1ڌ;6*El��=%�|v�i�zc8�P���j��rI��45�̩b�a@������!:{9��g�� v�{Uv���>3�D�J�7��s�y4�qb���T!ܬ�,H��h�'
�σI��KE�.���R���Gg�J6XY��zL����f�. {��2(y�$D�%U4�a�*`��[�a��~���04a�����d��nAǒ�b���S��&���fz�g+��ֈm�U	 F��m�M:�����m�(b�S��f��6ep��S���9��L2	]
$�T�%0B8ǙB/o�4�p�dreI�mǌ��_�5=���O��	y������:���75�� L�U�����Y	A���=vؕoq!���^�$�^ ox��oK�D��.�E�GZ�F�:+�+iߟ��ޜ��	�\�CR� ��T���7H��7Eh�cs�7������6��2h�3L�^X��,�����m�66D���%v���3����Ddv/����Kp��0�}��Ts2M��rcA�ᙡ�s�Jh?r9CI@� �6t�1��d�p�'o<,׀'8�^Pz6�����9�Ԭ��@Q|X~���`}@Z���_�<��	7(Eȸ)&A���/�}r���Q)���lH���x��u�}��t�N Q��Q��U���ؖ���t�c"Ƕ���l�����#'|,p��h��?���N���*l(I^�v�f;��~� �Jh�����%he��r�
�D{(P;r��<��UiS:����2���ZO}�9�Ǖv)��`���z��5a��39^��|�+4y�Fg�1LO�y���b�E��/�M�r6�G����ѽ���UM��C9��wV��%��M�L������cB1E#�<�h���Z� �����n����a�	�,����E*����pJ$���9���iԆl
���%��.fnE�'�)�m)m3���*�.�(��h���*��h���Z����&��A�쿈HY-ӼhIC�j9��q�2�˒�Kx��
x=��^]��A�V���$��у�)��g!�dn�?��hW
�1$�I�z�ڬ���>dk��d�&�^2����B����
gt�]�6yG��d;.(�C��nۈ2�2�d�s�z+����Klp�W&*�{,s�����?�桪� tH̴�qn�g�'�!��2DNU�R�<�,�M��$�������;G=�wb�{x�[\}_�+=4�N4�u���&j��ۣ����U���'޴X�7���"�>B����lI9��A*�����R�I�3���L��m���m��Sؤ�-��G��$ox���g����W��Z�����#Y���Y�{�p3)q�̳K�o*ܶ���.*@� ]Z�}��M�l��줡�-y�n���f�H��ad���{
�|��Ғ�@-11��Y� P�=�H+T9j�^2�
�D�(��D����h�Qf�P�+B��q��m���N�zc� ��������~	=�|<������2�Ԓ�?h;ϟ��M^�Ѻ��`�n�H�� "d�9[�t&8YE�o}�!#j�axN�Y��BG��tQ��^�ȱ_����oI��S��wMB��8�Ĝ���+��Ob�Ί'�[�|�t��j�tY�"�V�f�j� �2ǭ�b�Tu5�(1�c������i�U&��h��k�'9�dQA�oj4�GÏ�u�o��(�/��Σ�q.5_��GʚÿE��d:�� ����P���[����V��G��d���`���]i9�G�(�@'I����kA�����Gۘףh˽Ec�0�Z�$T<^��y�3�)-Z{R�7
�c,΀.w�NR�2<1�\]�S���үY�k9��1�0&2�G�/��G�!�	�ڇc��F(g���B@��N���%������� ��w�SRU�E?�pq��J.Ξ��I�9s�s��:�Ɵ��7t�sc��ƴ,��^
�to�yS��v���VԴV5�EӘ*�� N�T�@��Y<�O�ٮ�|�|��)��yh�uY-�9Y�3���CǸ���Z���e���0h��.j�~�������7�IĂ���I�݇���m��͜��>��`G϶��5��+���4hm%��n��2,��i��bM��He;��S�-	�r0��>��.���>pDT 9�5f��=�#��甦�ߩ����?��Mu^�;{���O�S>�`q�;�-aG^��{�}��'�tޛE�%˱�@� Ը~�����^N��!X�4��<5�Ny��ϸ�O�N�VO���=4_�`�x�q7i�k��t��ʺ�1�'���ąyղ���㴀�� M�#D���b�&����spb%=�2�g�k��"ϊ)h�AE^z ��mw��1.;��B�["0����Y�/MNT��)���䋂c���=a��9>���}$���g���~��f�R|C}�|�2#7�0>�]����Z끘�:�e�^ԅ<��V����C�@=��\b3��xE��`���(��h1�t���9
�3��تY�<ީÄh_��;�� �*�\�sS��o���M��^W�E,T�� Z���A'�:ǆ̸&�}aڜ�=�q�Ճ038���9��T�,�֬Z�i3�.���^��Z�e�冄h�ub^*��a`�����/�\ey��1��k�������
��ё�0�g���G����B^�u��?g����@!S�ZN>������tO����UJ�U�xz��r�K-iA�n����l�OϷb�����`���(?(��AJ����4�(e)�*��&Ij�n��@�`lt�^�n�L{܆�4���,ļ��Y��������,�Tr��h��G�r��_q�t{�8�����C<���I��J4�0��ӣ�+A���U�YٔUK���i��i�c�/ �ʷ�˫w-��n�T���G�֘����\_M�EE����i��;s��s~:1���glmܶ�GΑ�'W�{��=��Z�gJ��EtJ"q�rq�G��S�EPE����'�K�u��@Hp:}a��_zmG#�s�G��kZs�/A�E3�?urb
�Ysq�g��������0�Ž
fP�����5���	]�tcy<�<Z���yֽ�~���b�<�9��]�����cZ)ӎ62w��`�P�j��s�]�G��+���k�7��*H9q�|��f4#C���qb���E�֠��Þ����:sC~R$(�e�9�P=�% �5p��.�>���:lW�!_kO`�&�pq���.c��sd@�u9�/ѾM�#���}��k�E���zvӐ��\9S�H7��d��#?Bz�'i��:	a��/{`�?�_,cG�2�����:Y.h/f.���":Xq��މlm?���Ǌe�eG��m�,Bdg�p+[��%���9��z�#���Q�H��3R|Ra%�V`���́Zl��/?�����I+l�Oanؖ¯�@�'5l)[�i��k%����`Z(A'�{�HSR��4�7������W������=�TަR[�7�z����h�U���pyfN/�O�� l�[+�_Ȕ]���v?�0-������몭��hF3�#�"��.�{z4D�9��-5�oA�k\+!!/F��/�3(6BA��74oo�J=���{��sZ��p�?(�mr;�d,�R�F����n��G����U���֩T �8O4Q��'�否 ���H��	�V�l�\�#���+l���_�#Fq3�%�����p��x��v�~���T�Y�k� J���x�Y�?��WѢ����a>n|��0{	Or0�NZx6�eϥ(�E	1)��yoEw��Ny�@��or���:���hsn$y��hfa7!�uw%��i�;͖stF��ª�CSTA<C�x4dO�6��*�Q��E�2��7��>��3���|�"?}K?t��
&nC��%y���x)^��%	:��Zݩ���z��Mo����e���T0m~v1CN�&��Mu+��TՅ�f��l���3�G�凇�������Ϥ�G��1	��Oxԛh���Q�Z�ˍ����m�F[.[�	��E���J�^��Q�ل:�a�`���"y�%a]���ކ�67��c?�X�<akdm�O�E�0�ST3"���n�'։mL{�+����Ok��<50$���PX��� 2��u��~�-<_K��y=8!���"T��6&?.."G���Ka����O�&�M�4�LT�򂛱��4��_o�<��	�O3��Z�e6����e w�2���ڜ	
�W���@7�&��Uз��G1��&�;��֛<}���|���P���r-�Q�l�2����hi�`���3��e�_���hժ�5ι~M'�Z�l(y���������.�Ds�5ZC�i��*D�ﳈ��.�q�
����K
pE�==�l���1 [3�M����1���| �֥A��]SՖ���u����k͕!Hw����M �nV6��c�+�&|0�m�	�=���j)��]ޓ<Ǎ�ַ�s	�+o�4.�p˷��,��"= ��4����gK�<�O��G�߿m�nQ)6d�kY�ބ�l%�#k���&�ڈ���kkW6)��/䲿;
$��!7JVGo���K[����wf���@�4�+���U1L��@/ʂns�Y:j��W,�T�g��<�%�lT��=H���1�o{͌;663�J��4�:��g�/���>p���h�Od�?P��@�-�����М����TFw���c � rG,A�����as�\LʗΝZ�a�LH�]���O���u��@�O��Ո��rC]��/�O%��V:��qzǭ���4�T����(2������D���nss��	Bk��ӷ������*�m+������$�M�M��A��\V���9�2��UOku꺛+~���a���Iݱ���dZrDf��fi�%�|��c'��
���C��ܭ*'�������luu�:F�T
�ќ�bM�yd�v�2V��&�(�7��f�Fl�+�19��������s�o��ѧc�����:���K���}�C�ô�-g^�A�M7�w�0�����l�O�>�&.3,�eLލs�nu��d�{!�H���&�	ذV�ŝ�3�)�3.N?�rJ��j!ƅ7%�"�ƩQ?�FC')�f��{$sb�Ȝ��d�EtE�2�F5��8-b�F���~�]���$�;���y� )ɣ���}޺�H�C�R��|�������ez3���N}�cA|)�{i �s�ƭ*�W�¤�F��>��Y�΋��>,��LIäKB�fVѼ�d6n��}=.���&;��M�9�z�n^,�Fk�!
M3Dv��>���ݶ��puHW�8��#J��3�.��}����	��0�Y���;��m�c��bj���*R����Q���{rx)
S���Y�����
��������՝N�f�l�_oJ���kP�:&F��*� �k����Y�0�F�s�A0A����$w�����(;��P�3^.F!/�cU8{�ÊQ��ц�Qz_=Jl��&�2�%ZDi!�i�����S�[E �V�����O3_�^p� ��5�j����e�x�;]6�eT���pPH����~{���msvό��,p'���ʡ��l�b�C�a��|2�nu����#{�oH�9���YBR���֔W�J�ZYʳ*^�8���US�0=��Q��*&�>��˺wߠ�b�ڿ%��;��WS�Oڤ�[
p�k!�k�(�c1�џ�p�9�g�\ŏ�`}b ���J[�5e,����0M�L��r��@5� |��q ;� ^��!��̙��agQ��	m~1y����T�ɼ]f�l!�úg�+~���Ԥfj�^�
ߋh9O�|)���]ӷ�$=��k�l����ܴ[�H�֒9\*=OCQ}���V"��6��k$��#5�A��b�t_����������J�Ⳛ��J Qrɛ EG��K��KK=��R�vV�$��8�`��7�Ra��{L���=�u��0�at��?��k�Xu������V*�Q�L�Eia�������<��j2{�Ft<,�
�kX����p�[�x��b<����q��̍k�mɞ��j�P����+r�?]�#>(�$���6��)��P�lI�^ʔ/��c[rd�z����&p+ϔ��p�{Ϳ���<�
_��50�Xj�GH}���՗+�����b������hAO�MQ惺g{�����)�>���L��[��q暺��2��A�}�e����L�T!�P�1��3
2���E�iZ�k���E�� ~��A=;]���w$lD_��~�y�X�}���Np�'��Q�i��N˽X3���u���''gH�����;��'��b�bP9M��k�2�e�Z4�M�s�"��zm��胖M��|i����>L��-x.��kl@����;|�ܰ#���G���8H<de�#�8��N�a��J����WQ����I���&��`0g��gA&��b����y'e�GϥDG6��H<�H��Dm8���	.C��_e�f�[�퍁����I-�V~ѵ9�G|g�E���=�^��mUy��f��45�M#�����14�p�H��lFQu�Fp_ֵvuC}:d���u����0�y���X��BN���G+����/�����m<)4�AzOɢr��&]+c����[�=��W�$KI�j��e�}s\�=QP~�u?���h� �Ax�V�����4#P����w#_:���J��t�ڴ�ٜ���T�ʷ6z���2g` ț�5:^�"��Dꤾ=]���uZx�{uC�7���Z��� ��E>B4�!'���X�(���!���D���a�gBT:��|}^l$�����]`�;��-끿��c���~��,�
ϔ���%�
��Q�m(��6}����AɆ��h������$�pԷ���97����Ƌ�~�=6�P�^�WY�h�<�����o?�AoS��{�r�FN��a�AE!"@":�.���a��g�s���J�V�]�w�W1���C.�ycf��OQ�ئ�Tyj�]��k��ۑ��Ow�A^❽<��/Ɋp+9o}��V��M�$c�sv����=k����WgG�W��&�)�"[���Lw֛X,B׶*C�|;vH2�{�ܷ��܋nx��nUQ�Ar;bך���ؑ��g�YA�R�g#�Z�<[n&��-ӂ<��E�҅k?sY�IV*�������6���u�ޚ���(�e�ao�*Ȧ�)���kJ�BK�L[Џ�LI`�ow�khm<Ϊ��`!�I�W�P&!�3G��:��]U⠟��1|�� 5��U�Ò�8��e/TګkZ�+0�|Ƈ�q�ч��E���B|9�(�e)��lC~��x�&;Fл�(�n����r?�9W���(��YV�tWh�!C,H�K���\H���Xg��� ��������ܗc�� %OGaԱ\(�e3S#��O�/�4��-���B΅�;�j���6f�G3ޣ>��7/��Lz�Ԙ��-OT�U~�,ك}f�+�7�����������d���C��NھC爣�����E�j�L�gR�s�̤A����6�އU)�~J˼I���64�H]ߢ�8�a�&nW;1�x������l�>��qD��,�6�5��7::�H�� ���ӥ�iw��q�Q�$X��=����V�cV�;s �D��l��StL�2ĺ�j�^���'��XE��M��DNI2*����v�Bg��G�q����	9�<m�;|ɠ�zR3�3:氵�ܽ=�������-���k]���&��*ถ!F����#< ��5���������7��AW�Y��L�e'}�3�(�����s
��o&5XS�3�f�
E�xĄ�aJ�����?C�WH&��,l�(�N�`��Ǹ�_����4 �eG��G����O%�ڽ
~�k�S�����'s8�|��dv[}��V@y<4Q�z�X��r]CI�-M��>Z��~]`����JvM0�0�{���f����|���Z�o�7W�u�\��[8��!�?�b� ����ȃ�����Ahx�+��HE�Gޭ��wA��܄	�,���@-{�~g:d)��Qx[[�#�B���r���B��K�N��rߐa��d�pa�t�I�8������G�������э�f�]��y�����)�94pד��^b���x������ק�mЕ��{�Wf3�a��p�"��_4�qȀ%��������c�������U�͌�Dvk:��,��p�H7!��V����f���g�Ot�&f��B��:=�(_�ܒ(��S�i��%H	9K�������nz��	�]�2��cp����oI�-���T.-�Nכ�#i��0���
���ѓ�kB�ؾ�~G�m��Q.�qzf.y�ǋ����	��V瓸��Os)^��Ղ���u�i2�b��k�ޕC��ҙ!To�K:��c��`��ba�����O+367�f�K���AU��W<E����9+�鏔:�h;}*�|L�:ݧN�m��6&/�������+��6�V��f����\P~�"H���r}���y�Zh{Y�W��~�U�5��9�ߌ��S"�1�ѡ| �LޥP[!j �&�S���s��H!�/ЎO�2S�WZXNc�'�2�EWa����`�Q���z�1C���ag�/��ƫ���Y]���N����Y�\_�/�,}�s'�v������p��9���j7k�N߽��'b�q�Oe�
�Y�.��ET7��xM\��5�b��tI�N�*\k�S!�H�J�Y���q&�R�7`øn��h"J#�QPű�tE�t
w�;�`	��O� %��H˥JiHb�w�u���oԱ���`E25]�ѝ�����W�umҏ�E�>Q�`�^*��{|����/m�KY�:ꝳ@��*f�J�ǡ�7b���޹LEѕ�[�3����e�������S%�h����;g�i��d�r4��Dj7aq�l����#��1)�_�^����}Z�3!a;��˽���&��gVKCI����������}H�AM���Ȑ�ǘ+
�=l$�$�����H;��/�1nNjb=�5�ܜ�5��O�&��c�p>4
ux�K�̳�}=!����N�{\ρ,L���܃�玭�`��&0��A�q�.^�R+���R�����G�h��kR<��Q��zE�NU�X&�|��%B	�T}��.V�/d�r9�	+qˈi�DU@��3m����%���Ps9�v�Ȯ��I*�t�D��HLU6��#?���\@(i�@��6GX�E�
������˩b��I[�G�$b��z��J2���/ͳ/�&�@�`�����O����J��A�"ˉ���^��J1�C�m��qh��r����F%d���*\q7��q��e��#�����W�1��봨���(���pÔ��������Y�}Z����S�u���O��A��c�=0�
v��f���Lz��y��F�j)�u�r��Ԟ�WOWh�ޱ?�P�G�Őgi�A3�����U���]g�}�WH����.\�3a�r0�:�i�����uj]C�@'�9��?� 5F���R'�럝a4����մ���X6������,|,[�C�
p��pQ��Z�����C4U��إn�j���K��&B��Ā�,��y'��lWy��U/�]d�p?zTMC����@��ụ��Ӄ�[��&��Qs�9��:�w�[c%W���H�I[x"V}8qQG��\D,ޝڡZ�ψ�2�{t�<̶�B�;CN��)�(�ry2�d����9�O�`�4*f���_�UӅy:����=��;�$.~$.���0�f��4�t1�VԞｊ}y�s��ʙ�X�۩'	%��=Cl��l��<�z�N�ҁ#0|W]����Q4����܃���p�lF��p�>�!٥��8�ǭ�I�� !Z��k�h﹒�7��Tfͣё����٫���̌�����)1�K,���52�   n/���~����F�)"��}��65�Z>dVR �A�%<^�>�!�������Uˊ @� ��:��y�����x�9��/:|Wxt�����\�ċ�>���]a��-���N�vG���⒎0�,����c��
��Nͯ'g/���L��Y)|V��8�DR����%7�P�MlK�
�)��1�=��7�1����.�ǔg������ý�����IQ�Ӡ�P��Ma��#~ ��"z8��pk�0I�No��0QF*�"����쟲 ��$�5Os�a�:,Ry�������o��-�~�S;��$�:A������吚y�r��K�9ݽ�Y��a9�M��4m1�/��X�D�"���	�i�����?�>��w����ހ��	�����np��G��f�9�T4E_���_h@�*KJhD�~�$��$���=uX��	~��u�n\NBi4���2ꙃ�ϣU�GԴf�z�W!�����@v�'L51d��<�xMޫRG�����:J�(F��q�_�ʷ���������KL���z�=QdJ�r������� ��H��~��u�)�u��L���\�%c�j����1nj�e����ju_���9�0{�ѐ�-Y|���Q 2���^	��V>,x����c�)���E=n��AQd�A�B��;F��x��ō��D��jl.�%ӗ�̱3�Y0��C�3�t�<�?�/�ڟ�����8]szY2�m2�o�������P�r����2�}C��R����� -�ЊO�pnx� lѹ~���{W�vH�>�4�\_���R��r�S�OA�tI� ���� �D����|F�|k����L̊&�����	u ;����{ˮ���2�Ġ��5���h�pS� W.H�R`�*?�����Rj�D������u�g�Y��Thx`��9��ԡAKz)�-vQgQiAk�wj{za�_I�H����iM�5R  �a���mg�͵<�b�Z�1�FGs��	F,����t�a����^�����hN��	���W�{�Nɝ)ep��N]�-�3�}�O�Ȉ���*��h�'�Y�3���Y{������dz�{w5��.zE�4��	4��yW1'��N��<�ꙇ0��,,��e&�=:=�Ղ;(X�FTc�ɏ�`�Sa�8U���N�c�W6r�J_ף	�o�6��ݏ��N6zb�YQ{
���rPċy�5���>H�)�j��z��{�pL0lR���6�_G��X�<�"��ai)��b���Fg2�S&ڂ-����l�3"�9J��,^����h6��$����*��v��$%YЁ2H���P�[�|lt=I�`�-����l���~�5�g|6	�%��A�K<�к��=���3e�cf��U��g�� Pk��G9�x��O�@~����b�#�"O�4�Y�������INo�d�Lj��\�[m�!�M��db�mЭa����Z������*�O�<�,a_��_ �2q�~	��3Eg��y�\����Ԕ��a�;s�u���s�I�=Z��B���
UCW�}1�~��T^ܕ�4#�f-0ַZ��r����p�T�>@�����<`��_UV~h�pBVS �Iq��A_
�S3��!uS���hQ�g��nh���"��M � uf�҇��#~`aC��$�)��9H���}�ˑ�.���di
i/�9!�ݦY�Q0P?_�nً�A�-�6�t���9�G�Ƀ��֦]��
���9P� nnv���>��(_Ƅ�������ӗ�}l�r�i�QV>�u�/��=,j$X�ϥ|=�l��t2��o�q���W�2�����>�J8�z�˝0�ަ��!>ﵶT@��^,�ߚ��r��Y�Y'��S�|�A��C .���csB�RHD��8������J��@�>�UF��/�����Xnᄒ�bi?�����R�$ۋ y���DK�uĩo����P���}��U!�}+�K�K�´Z���1S����q��|��,9��j-��<s�8�{��$��9�BvW�*+A�7ځb�Gq�J濷p��򻆕f�rH>�u�UC�"��_m
�^��-�s�aث��N ��aMZ\|�
��2�����M��_<N��;�v�/���J������T���Hz��B���I�*MFRe�{d�nc�!3�#ۣ5.K�;;-�	>��p̭�c_����曌t�k@) � ��5Wn�� �X��	�fcO��`O��=�����v���$W����T�wN�PG�8Ғ�'��ष��4�^H0aL>I���
$>*�<�DV������/�l������>j
�ў0#�4�`B�0*�9���k?�Z�6QQ�7M3a�����j����t�Oэȱ����H՚�*rq�4UF����z�>np�\�-��e� Q>�p��t�Wa�����r����S��o8�?n�1�2����F�ٓ�p��+*�oy���[�р�d.�T�]��>�ߛZ�^sw�\��0_d�U���gO�������)�?C͹������h�>E���W�u����xE����"�,Nd��z�s�������t����Qrpsy��9�&�-	j��-��� )�8�y}��8�ZB=�;�,�]��9���� �B�ჼ/���i J4κh���
򛢶2񴉲W��A���V�G��o�@$�c�'D���� Q��P���63`i'�[�UM�t6�0OEe��LK�����l��h�u�HUtc���E��۵������I'4�J߬�8�Dg程6���V���ޡj[��Q"�4�ߜ��`٘)d�Af׀t����"�'�/���T�#�<�->���Cdb�GE>ӈY�9�)�̈��o�+�熯B~����~����)��Q��d~�f���X[]3H����2>PQ��:�]HK"��㵞&�]G��k+<�|`a���	c<&�Qqf5'�Y��*����kҹ�]ۖ���	b�Ԁ^E�9R�9����:S.@ +�m��M��ۦ��e��X�IV�#3}h��?���
|IJ�ô���v��Di ��g�:թ�ԩ�)HaN݂��P�ܹ�^� �Dڍt�s��	l'����BY�7t9�=�N�Ccb��"����4�^{���;�����iNc\�rOүre�~#����&6���5e��ZG!�G���4U�Y��'�눷&W��jyI0�	��LQ�<���Aw�O�h�5H!�~.ʌ4b�]��K"g˂_���Ծ{v��H�)�V[��qĮ�QqH$�"cZ�M�R��Xc�@��P�2_`�V�,��D�����A��J'��xs��6r�s|d�D�J��r	�����
r>Y��>��y9T �v���	%q�L?�LC*AP�vA?h�=��	V7sOOaR�[�Jb=S��뚌_��W�]qn�T{��a������%�A��z/%�@�� F��d)� ����?�%�2j�Y�6�.t1ӱ+���x��qU4�Y����Q2�P��.�ې��