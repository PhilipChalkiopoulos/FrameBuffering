��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6� '�7mF��+�Q~y�[?(rЄ[��H�{���Zh�ƯD	C�o��M��+�I�J��]<At/E�8~�8Vp�Ef�'�ǫ��ZW� 	�,�*�Y�S�gF��ӏ��L�2��-�ű�p5.Ha���H�1���� ��h�ڗ�h�|7�F~�QNy���RŻuC��m�4#}�ND 4S1H ���J����Ě�XaȚ��.�}x�M�W�[�w�	Y7�65�Y��6�4S�D�c��sA��!�Z����BJFAϛGw���V~er��k#!�19'�^G��N8�9d�~U���3����R�be����w=�O�>�[��n��U=��Z_M�@�:%�� �y�{����he�������,}Z�a؈�_�y����e�I0"uz�<�`v�2�Ih�����aY�q��G��4U®�7���u�Ya�X���SLX�2ո�ol��Iٟ.�zSoF:,��۟3���Kq{���`��Zȡ`U��㊿M���o?6�ɍ�wp��q����f���������o|LI�E��L�(q8%8�ɦw8�aՃ��ÑP�Q���Rh5̒ �AP����P!�R%5�
�^d����T�#��$�/��##ݷ:6�=��+��[[i�ڕ-����oXc,����	Ѝ~��"�'t��G.`���Ru�_�I%��܎<��;�?(���:�>��de�3���w��E��hg�\�D����M�g;��ϛ��OC��B�ÉNj�ƾZ	k{��7�BY|{?&��{N��GH+�};�)撋�]��N�p7!�&��
�w\Mڟ���D���Q�`���ʽ*R����=�<���`E f.�6֕��]�e
Y>x�a�Je/{��Ó񗄹c��L#�n���kԪ��%��6��A�x������11� ��'�?-h���N�B�hx�d�z�ؗ���EE�k*��"�KvV�b�3�����c7��U�Ӑb�F���İ�[T�c��)����)�F��wr����BH>(W��iZ���g�~��1� �X�%G������D����o���ң�&�s��[ ����������,Eg��^�$�'ù��V�~�?���3��S<C�0��~י�Hۛv[�r�ïcI+�;W��Ѕӂ;�?m0@
����ܯy&�L�xE��y�G|:���ְ��#D8N��|/�펾V��BQ����-
V�!_y`�
��JC�X�6��紸����r��wE@���.�:��(�~�^�>a�Q���^�Qm�
�y�{�潬�����*�{��A}�g%�����"��z�R�a�e ��w�ص��>��U�l���Ǳ�6��V�˜x39hO�B񰉅6�y�P�p��hW��Dv��2hh��M>1��26GH��w��,�)w����Dًt�����zy�~V˚`��R'�e�:)CF�}�T#Ro�F�����H]G�p�F(]!d}ߋ�a�m��ԟBȰ\�0.%ӓ/������t]�0>|	�8w��du0�4���h���1��)S��7��0�4i�us�/9A����跞�7�W�E�#�u��g�%k������ک u�ٛ����~�S*����k}�-&h������*������dO<��l���]�5�KzzEH�L"�ҧ�OtOoP����a$W�8zwxkH)�J���7쵛�����c��c����rC$j v������{��{���M��"n{��L��C�ʍy��ͽ�b_��?܀ٕy�*$�E�5ՓP}�����T��	M��Fi��t�`J�}�\5;�z��Y3���4�f�P"'�qx`�g������#�=o|���t�ߥ.�/8V
9��L�yK��U�.xB+ߦS#�E��y�"(T*��-���&,<H�!!��C������5J\��9?&�d�"I�>R��ޚ�2�K�E:9c��Lo,�w�!_�����t�c��G��M4���m����̾WYiX�h��I�_9����I��r�K�My��jЊ�MR��N=|�	�n2ي���J,�4����Wm��C�_��2�- kj ���V�&M,�K��nQ�ʐ��8�Ed,"�y[����d�����TѶ\���������ӅM������[u���8��8��X;�n4�`�'��D��������ia�+:��,6q�'��_�vלlr9[���/�a�֪{Ny�z�6� ��녒ld9�j�1�2�=(f��Ŀ/y��-ѭU2'qC@��!�Q��!����'�����d!�b�%?z�$p�����g[��W��axܕgCD�-�v1�gT,���X�˒�Q(�� L
Y(��z{��D����ΰ���sԻ�p�ϸ���-��^ܜ����7�lmI��
�$#Y��p�g���W=��4N������y�����:WH�Xz@���ܒ:�����������M�;)K�b�fn/��^�� �p L�iwj�HFhnl��"�!u $�����_�����ʉb���+U�:�鮍���۱QA��d��>����t���z��J�� ���z�1c�(R��F��!?�� ��3�8���_o?<�,JсQ,h�f��?��IF0�Q"KwX�Y�<P��Q�gO:Wx[Z3�R��t�p(��ox�P���� _'y�q.Q��OH=b��]O\��*ĭ@��uK�4g'��9�98KXd1�>�=-����*m[�Q3F�.���c��A���
�~#�͙ ��oc��H�>PzW0�:����N�Z�BO�9�T�iگ�WV7�?G�C}��VM&]��R��e7ȷdx�4ޏ��P�$R�G�wmaS��kN�[�J�t�fV1�h��x.�/�����ϵ?=O|(	�=�� 	��{D�*�~��,����>gІ`��
d�a��0W�6�pG7����z޻c�r�wb�n�����r����:�ؕ�h@��G�A� ��*�S�3b��	0��2��<��q�5��&�t�Ű3�H}����!Ze�ȡ�s�O�����>>L�O��|G?��dê@�S }��	��]�e>N9\8��i$s�Y&L�[�%O�s�<Y��SH�Ft��L���s����q�k)3���G�����g���2�)u�e%l ��?���䏺�H߀U=�*����(
<�R�F�LV�����$po��1%st3��t�m��%�,n��ڠܬ�ɭ*h4o�����/3�y�NeX���zD�	��ړԾ�g	(��Çq�f��}p4�)3�g�q. 	U� ��J�唀u����Ǧ����jV���U\�Q�R$ݿeY|��NX�� iZE$���Iz|�Y6n�
��$� ���^�W���PZ5����{�	���[4���Q��>�w�U�NNLxAQ KZ�&=�J,��(��4��Xn\S��Z���Vy�2L+�Qܫ�%g?�;��g�;�˧֫�?��"x��Z��8��բ����E���&k��U�H."�;/$�{hϏ�D��t U�%�`��Z��Ⱦ�<y��C�4�#������L�{{-x)_#EkkҢH!	�c��n!�̎�VD�e�!>�y��l�����3�[k�P��d�F�@'G��h.�6���p��%��I�>1�J�p^z��eW$C�&w>:?oo)��>s,V���G�6��
�x����Ĭ�|�+�u��,.�c����г���#lw�v��Vj
UdY>�o	g����N@CBd��Z�uSv�]�����qЋɏ1a�g�*�)XG6���/�j{.&���B�-,�5U���g˱�	�c�ǑA�i���E���TT���C̱���ƺ4��U�A0�c;��ʷ�@CO�=�����Nrw�'!_��U ���ȷ������X�j+�m_ҳ)d��E��J��1�6R�*A��Qr3	�O�g�eK������s��@q:U��.o<`� ���r�~�:���Jo{<�t0�?���X�v@�R0b�Gp(&�­����K��=&��?%q{|�y����O�>�N����m�������Y��Ţg��Q��0#�^E�k�	��nLmJhg;��jM�\Y�]J��N��q��,�(���]m�P��'���nr��i��Lc.���tI�cf1��Je�/�����(�L���I�h�?݃,h�a����o��8��i�.,o�p�J�\[�pA�q��v��"*w�cb�'���������?�'P���i*6�nwz�?��z����fR���*ĿLHp#�F��ԃpf���'���#��i%�B��3)d�ң:�0<;P,�	
[y�_Ĉ�V��f_�߻�r��K~�����?������ ����SP�t�{�K���'H<Z�|?I��/�c�%�+��I	���q��Jdc����ٺ������e���oP,��_Ihaɨ>1W��?k)��&���N�\|H5�q�������;��
�K��_�x�^�/gŻ�
_����1��Y��_xit��ȥ踢#ݮ_(�l,0b��n�bG�L���/�e��Ӗ�<BB�]a�b(�aǮ#��q.�mׅ��/uC6�����Z�V�����Z�gtgM���l�E5|�����F:��ժ�s!u�eZ�!�}�����aM6�o�ن}q��R��
}HQ�<g�&�)��yÁ2�on�v6�{���d/��b=���d�]1"��Z 3`��|T�(d���r��u��33�?����� oz����3P��7+�U��|o|&�S�d�M��s�S ����Cc�hq�Q���?�x����EM]���{|�7�=�����%YNjq������c񰺈B�\4Րw����%����`L~�y�������?��ʦ�S��)T��u?$�c"i�t �|�߸*��Y��B�k�����:�tE]��I����E��橿��Y!cS�D� v��o� �4�CY�?C;#������ּ����q>��I��q���U��?ֺ�?&w��v���R��d{��h��{�o��;�'�}�|�C��.ق7�#��0����&tyf=����[����f��ۗ�]a/��H��;8&t�HVWOj/��ǇAE,n[�ko2P5��K��-g{�B ��󟝬8�J� �mz�3��\�0z[.��{�Ðq!�>*��W%I���*o3㔋�4���eW_�qH0�6�v1���d�t�`-l�d�؛�jli�>l�7��Vպ^Բ���
�l��1��'�1��B euB\��׌-a'��6�8(�R_�������P���"@r_�C5x�db�z?NY�i,@$���`�Wۖ�[�IyĐ &�'��#�}�	U�S3����Ek�,c���ڱ7󠕀��$�N�|��� FZ#m|
�D��J���aׇ�8��Q��k"�#���������N��!�A4m��_txr�?'��hB��3ǲ�u4���zrL�a�:s��෰��f���kQ�?�j�>Z\+ob+;�����I�T)@Q�x�y�wT��P� 4�a��!�#E�1V���e`,'S��I�
�x���"����+M���Y�4��n
^�Oj\��vF��t��]�����aJ��[+$�o%!L�ۙ2`U���k���T��?�Gԭ��jh~�N�+$y8�B./W�,3���?�K尀}M���MW�mE.>]&W�D��F��4P���'%9�b����t�o�p�������3�ƨ�]bQ���M����2˭���G|��J9��B��E�8P��R)��cM�إ��ޙ>YƘP(�:D�{Y_���~&.Xx�8��Y<��IsK$�V�i������r!�}a��q�0��왡��9�n�'�t�~^����C' oU�眙�T�	��:����"^<�+��P��Hx�V3�,�
��������M���Q�	U��O����
�So��� !�SK1p�����h&fxNX�_�y�#�?j�V��+��'�t_~Yj��b��g��j�غ�d&]X\S�7����\�ޫ��O���7qJ�п�,�"O��σ�k�̖�\`0/E4�k,�&�x�T�)͋��h6�C����TEV�(���/�f �u53��Aģ���{k���Y��`�r��'��K��3������b�����	�1�0�u��n��z�2��h����X�^V�U�y9L�̦�ZL����r,��yOY���lrO(l>?�<�&��w$�}
��2S��?xݜ�Ib��1���
).�b��<O�é��	=i�s��%e�����ݥ,�C�o|֔��,{E$�t�|�x�*���.dl����EF{>4�%���Vp�,ka��0�=�c-�16W�]��#������-d�;����O��=���;o�WO5���:�x� 6��]�y�ׄ���r��n�!f�
��oC�;Z�CE��h��uM,�?}�qt�0���k�Ր���А��A�|��=�q���K[.i67Mpgs�~�_�E�ֿT$n���)����L�O��w+4(�8��Lfyɘ6\��I]����4��G>.�f�쮘��܋p�x�j��}����K��݈��Š���v^�C��<3�C��u�KSf�Mqg�tLn�}̄����c
�{�'�i�$%U��	A�
�3�kM)�ݧ�08 
ba#��TZ�rզ�J�p�e%C�fIY��W����,�����]^jੴ��DW�#�IhT3o�3�v�ZYv�9�d�#�y~g������m9cpỲ�J�p���a��(�;�������阮T��]�W-���e��}�q�׻V3�7��UR���S�g�-���۲��j�%c5<������ԭ9�:�M�*���0s*m������Z#E�/������}��xl?Ih�4t��3�bZk̕B|��>sd�K�n�T�v�jٷ�Y����+���A6%�і �M�4�:lmlgC酮�T���؇�K2�v���C�l�����0v�s�nH��GRT��d0#���mֺ��	$�*8��~��
����T�9����}�����8��#�V��R�z ���-ְ�;!�p��j�ɮ$��/�"��;�H�슼%�7h`3��q�_'vh,7�o�03\+t�6-��//|���%Y��皒���.��Qd�0/���1;��IC�d^��)J"c旄(b��ܒ�OnG(��o��Y��Ȼ1��� h��ܑ1�g���_�R�(�������4$\�u򈝠�)���i�u������nq���"���P$��Ș�6��=�`Z����"�NjԢs�`e���f4�Ҷ�D�^Z�R�C93�
����S�vx�!����� ���̥/���s�cEQfj��.���Z즐�_����JV}��QJ�p)����g�����;j�s>�H	����.�O���Z�s��z��=��j��Cv�����<���e��Ġ�|£��/�7*YJeǜmŶ��I\w�OΕ�fd!�C���N���MŸ�w���d���"��|&ٿ��k^ǜ���G\43 �k-Ky�i���@@�"{���mbX'���i��m�]l(�ѦfU��3�}�S鞗"u������T)5�!��h����Gf�=h�|n��=��U�7�P{�vsb�>� ,����C�~������a�tV����=]�]��@)�I;f������!���aw|S'�[��T�Y��J�Q�"&��@˵�9'���xog?)k��gf�$�~��<�5���G��D��gz^�za�0E�m|����Uٌt/W㩒��]�c���'ߘ�� dL��u�l���|��x�+4���F���f&=�@�*x&��j �{b��i	�qf�9uR�����T������������.���\T\�Jg-h�Y��DB$:I�r!7#�걯1��`��%UZT��qjN�x���]1�ͦ+��f�W�7n^�z�x����`��{5��'<h�4������1��	�]3f�ET�C�ԛ�Ą�%[�0f��®�=��f=y���:�f8�R�ɸ�����̷��D��]�`�w��s��:=].�uy	\��;�$l_1�%��Y�	/u��eʳ(L��*-��Ջ��!�d�@l�	�F\2���"� ���`D8t��^C%݄�V�\�$�=�wvTsF�c�SR�-�
�x~���(��Q(+�%[�R���v�Gʤ��(EO��n����+�O��G��&�Tb�s��	(f�����g��#F�Fe7�N6��)kڜן ��mT'�ݑ�������� �40V��!C��
q2M�ޗ2O&��D_!Ƽ�#-�r`*؀Bwa'�>K�O��$D���<e?8�����y|PyỢe6K�g�5������Y�	b�K��C�ejk���V�V�@��ۋ������;�J�����aP�#%_�gp�-�i�c�n�ç��H孚<~eR�h��;l��1�z3�i�B�`_:���E¥��W�gG��]��,�x�(d����3f�s����h���U�]��Vq���;(��?�*Od�Ol�,��kCFz�ȿ.�F�>�o]
��N��?����r�>$�wB��f%�_ [Bs�0p�b&bQ4�I���hV&�ψ�:/��6l��>�s7~�"l�mX��g��:,	��'a��˴�2�-L^uC�3��l��`�E���/K�R6�}*��+��H8���8&,��%B�`�smϷ
�`�~ԻLݮ%�h�g�5$a��Č4,܄WQ_i���lϦ��0��AG�<r|f�F�6����H�
G[?*{��Ѩ��{.�����.F%&�9v\���bc���KIB;�}�Kt9��l>�Np�ut��w�6��u�l�!˥+��U*JH���~����"��CFЂ�u�i/�}@|�J�ېǽ`W�pD�R	��A��Z�PS���IE��I�k�Q�=�ς�#�l�#L���z$[���،����̅rL\�d�JS)�e��Z{�� �7��Mꠚ�M�����]Lt 8�yK$�"��RbNycV�41(�	hF	L	Of�Uʳ����+0]C��ޠ���,��{I�#d���۳�=�_�
uKg	��h!��7����70�j�C�q��J�nb�J�MCRە��:-7�Aՙ`�ö�Yt�a�Dt��G Y���.b�nLʒj}*�����UJ����:�����8L�~�eI�VpD1�rN�F�F=��,��+q�!\��~�*��|�8�aħT�Po
h�&Ȩ&��VFu"�w�LM�Ԋ�ќ�A�f���<�_ΪAs-�k�<�d�ghֳ\�P�(�t\�8�[���l����A$��nJ��1VV��(:&dSr+��5gw4^��Fk�A
kx̨�r��I�(jP�l�g8#Y��fd��s�����G�R�ŀ��O%���@}d$�^#�zc���RR�=�sL'��6�$��mQ�-�u �3�kK��b�x����-9�2���kQ��@T7.����0%l��|�z�҃�J3x�`<�g]o���(��C�k�_���{�`�3�m�SOPE�|�=��Q�
��A�b!��\�0�����p���5~�V�����o�K3�1'�٫FSS_�<�O^~欮pȾ��&����F�`9��"O�G�����*�@�x�*0!q�>ץA�gs���A�<m�>A(�A}VM��_���*���ʈ0�9M�ua'E����r���%-O���+�����Ab͍OɃn�kKW ��e�<�!<˩�j�g���F��簏������� ��er���#�f;b����kK�N`���h�H�fvz2� �1�Eʦu��U7��f��FB����t���(�O����K[)�k\Wpܡu�@U~�S �đ�W�X"��0��]D~;�����h�]|s��
]�f((�4|>��	ʚ	&�]q��qjl�a�������!#�)�<A���Z$�����~�51��ЭL��09����$��Ԕ)KC�?����'}��
�#C>�=�ެ�/�Y���B\��,��'��3�n
��݅����+}����.��$�}���l=��2)]z�g�}�����@9���<^��I�};��$9��N�h0��@��P��,�?X^F�fG8ayW�(�X8�NYP��G9�翷
7Sx7��Wk�u��2�H=�H��+���[o�!d��+hඵ�V�2��E����������kE\`M�a�biu3t>���c�Y:*p|�J�A��.fF����4Jr���K�#� �9�_�c'p�LY�R�g�������UC3
Xk�N+�Yyg��(��q���x7��WXȏ�L� |�2£[���Bؐ�<^��<34(Ѩ&��� ��;;�x+�װ��;��f�����
���������o s�+X�DY'����h�Mj���hF2N	#�<g��fVb�EDw�b�)R�[[�P|u�@����r.�#�[
n���"�2K(���]�LF�Tn��䈕���5T��∶E[J5���K�m�	�w+ani&*G��b�=gfN(���$�8�Dg݂~YR6O
	ץ9(9��FZk̈qhn��o���|�%��˷��*N�y{	0s	�5@�L��!j��J?���"w��Gc�X�o�c�8��6���~L�6�Z���� 
�m"1ɡ��ϮO��>K�x����m��rչ7Yu��m�*n+��s*����i>����+� ��d0��B���(��N|�u5�^�JQ]W��W�k�F����������֟lf���2�85E\Յ�5Q��D�7t���2�{d�\X|�^�`�U�f�/��g�����A*�1E;�H���V���1�UPi;F5/��?���#A��K�'-b�ߦ���5=+B���="�QC>�$DP��y"����[Ql��~}v�$&o�	���\���D�ơ�'���u���*�d ���r?�(�iLq�h����1D���=n�;�|�/>����&{�
�eV�䧍�1e% /:.����ˈ?P	��Xz��
��S����/>u�u*�ޤI�e���0N)a.����Yw�l���Gɉ4�r�c�|��_��ȅ���rEA��
.p|H���e������P9�F���n��F`���\\ \��W[������*tPx�/����㹿zgON���A. )��|��<@#0qZ��=��&���P��Z��?51���;{��
Ў��f<Хŕ:�OLܠ�I���<_̺4t���|ϻ�%��}���Pe}�9�z`��"�,��]�3.�h�.t5z�ʺ��nk����b���7�*�s������dZ�H�4�;�ZL�7n&,�-8\��@�E><�[|![�_Kj�m!����c�K �F2����:TX~ؖ�D���b��)�B'�`z�&Q�RcOj��-��ٽ�d���VW2�k��݊4�pgF���X�d�;%Z��'͐����V�+Z>HrE��hhc�`	�;B#���I<o���F��,A�ف���@��HYh,#��#�.se���N��s�>����GdӮ��85Zw�o7����x�5����)�O�+wFDC�6��uU�f�e� 
��Ip��(�����	�EK2X��aE ��+��~�u��݀n]��Amh��M�§,K��?��N^L��J�S���N7�B�m�G�L;�Q�l2��?�S��i�2�8�:�[8|�y��o�i���}��J`Lֺ��� ���Ǟt���;q����m)�JF�gC �Zz��)��إ����S�����1��X8�9`�H�r�i�%�ִ����Êi����'a�wmq�H�����~ƹd�5��B6�Ws��oR,E�Xo�R3�T��t�,42���XD,t�4�����Uh M�U�BG
MP��:�`��a�f;9T),�y�W�z��pZ#�jOT����ʢ�o��A��p�;�5��^$=�?�����1!2�N�]h(�oUŘ�ܦʓFT�������+v�m�ˍ�9^$?ip�L�s`�wC�A�P�va�U�9t�V-��ġ��1PĄ"bˆ&�fU�X*Z�Ѓg�0�Ȃ�����*GUD�hK�B�N�ʎM�(�$��jD'���G:������ſ]e���3�y0������t�<���x
�-����ruٕb�0�2�bB�ߕ趀���u�/A�\�ڲ�S����L
_����9>,l!�0���۬�"x�mY�e_r��Y�h��S��c�q��x�܉l�ACm��n���  y�� g��eӿ�#I�ߩ��k�0 �+�H�_��.l�.�e��P
z�7�73K5�sw&!�U1��6���k�!�W���Fa*`N�O���<,�SV�����������(�{M'tyc��2ڨ*1�8L	�	GO�E��5}�>9�W�^4}��:����:pn��sk
}x$�9Y�b{�)G�R��w޾;r��JGU����z����
�A�$Ӹ��&���rh�`��82񲙢����1���;.�{��;,u= J�z3�n&���YnBڜ�d��&j�}M69���{��T�L�~�aWc��Ј�E�Z�O�ǂ�s��_o
�Zw��-�Y�yZe>�^�b�h$���w�o���- �;�m��sw�hv��E�~�F8r�w. n<�;��r�E[)h#GӟO�@22���?�I=T���g<W���H{&���x���]"�z��CO2�����!�y
Γ�:)$�T�y1����,�>^��ɍ�T��� -�$w;\���+���p,e	����z�/7.FYU�ȧ���p���ᘵ��s h5�,�?����o_N��Y��O��N���op���z�}��%���)��B�`v����f�;=�M��W�����V���yߌ��ʉpX�"�4+V��l�[R�=� t�S�}�`)�����{�E�d�v+��	�=��������~�2��"es��'2��?�����!�4�o�Gγ��:�5S��i���q_*���~3�1�.��(#v��I�U.��#vIU��;![8&տ�8�7�6l�i@`����{����4���k�.rW�%�w�o^�a��X9��;8@�-��\,�ؔ'�'���*v�a >ϡ�5��N��_����fr��M8�ȚF���YͷO2��`�SA������L.��W:�n�P����E���h�����pK�ǙЁ%u���W5�����N���܉'� �B�$�|��� 	XP���$�lQ�8�9k��mPC�^ߖ�D�
�4��+�sXL:)O���n�6,Of�y��ŁД7���J���RHVg}Æu�thJ�U�ʕ����ʹ�R�f���s�M��4��?30��|h���7Ǔ�|��r�8�Q2�OgZ8���9��yp�c�q*|��w�>�W���]����]��VJ�X����M�����K�����h�q�&�=�
�����sΜ�'7�#p�Z���Q�P�v��*�Zk-�n�
�������v�ȥ_#�",á@�oP
�JR��T:� &@���+4���'��H�����-g,���L�~W��4�o���Eȵw�;����O::S����U����Hl�x3����[f��3	Z���n=����w��1v?��͗Y5�)�QΙt�ѹ�t�&����ɨk�w��K�־��0�$�hH���0�
8aUh�q=Y�O w�F9�\�>�^����*5��+n���V'>�tC��i��g�y(0�HS�i �!�wH�M���{����,H;��=�u���g4Y�EpK�RYҮ�Ⱦ���*<LZ�^V�X��/���#Ip�*k��o��AJ�N��ރiAtZ#On�m����ߛ�.)N�)� ���c��@�vr5+��i��L�i!�	�6�n����eU��Y]���ά-`.©x�J3�����ǰ7y�'�̔���en�P@���0��(���ٴnx�m5B�p�Q���x)r�~(���cB	>o�U��ZF�2�q�4�`u����M�{V���]�L5L�&J�yW��ŅN(|������� �EC���X:�H�ؽ_N� ��5A�5����aޑy��8骪N�]�z���tq�[����	����hsi����ܴ
����jLu�]�*�LSK�2v�N��s=T��F���sZ��ipT�ofdj��F�yGR%���5�>M-�������X�|�r��%�!_%�z*��	�|x�at-[��r�(r*͘G��B �NRF�m�_��6�R�ߔ�7"8b*�c�0?Y�G���2¯ ���+�ٍ�����b|a�m�oG��xm4MU��%慥�HT]<���X���ʐ*p�)'ϫ�39���E0��R&=���(����)��+�f���xZ�����|�ӡ�{��7C�+2%Ӥ������[�pe���6�r�9%�k��z�AUq�S,�l�@_ڟ9dXK����1��ʑV�$�5ھ��`K#�|;�z��U��2�cߝ<_���9"�?�è5e�͞��ø�]��� Ks8��6��M��[��iߙl�J�WN��:5*��5밮2�g
�0ӳZ�fP���Jt������J�s�
æ�1 �,M�i eA[���ǯ��Մ��3��m�ѫp�!�|Ε�%0�2�ToX�CW�?=#
��|}�c�e����n����̠N	%��i�v��/(���s�V�{��w#����E?�!'t������� �Z�^!��c��l��$0"�-����˖t8x>�	Li�!��z��)�}������ӷc)<�6 G���wE�/�� Em�]i	�"6�?�k�̈O}�ȳ�Z9S_:���s��y����K�v���oe���m���L���01��J�����:�-�0-��@�7@m	��uC3d!��ch��z\g�m�L����j�
c\�������Ng̯�UfP5�>�ˌ�W�;U��x3�g" J:����<�[�Sa��Z�9�z��H���q���s�+R�͖���KH����ƌ����M9F���:�:Ca?о����pi�,o�si�7XX�֓4��)-�˙7��-��W �w��@������:C���*65��X�\Dr� ��W������0�޻D��;� 7+Sl�L��LbHdlNA��ܝUQ#B{Þ����z�����1u��q�/����N��X��,w���`�����N�u0`����k���I��J�1ju;����G���ٰs9�#�^�G�ǋ�����M�ez�?�X�*ƋZfWJ*_�����{� r(=��A"d�ټ�1�.�D���?���b��I���UD\�����g�%c�z�љD�?e��\����BƏ�X��L�l��{���d.��o�4Th���/��&�U�&͚���͜S���@�9���ʤ#��L�����,KzV_�9"8�RϺ�H�Z� Bk�v�-��3�%�m�=�F{��}Z��ա����]��V�#�go/�e>���ךJN��p� �o^���H*�m%��/ne���4R�"g�;�˷���m�I<J�Ņ�1�R~��X��f�h9���EY�g�/�}����Q�q�3G�~il)��.��pX��\���a�j炙�z����:�E���9������SID�����ԧ�u��)�� '��"�1"�4�у���{F��S6��S��[��y��{l�j��f�s�uw>)R�}#`�)����+���I��N�j�Ba�5���?��������M+��y�Yб��Q3aɑho���I)�hV<ݞ8���h�PxR� ��\آwb�3����WX��w�]$.s:��[3�n=kz��0b�rE�{)�6��NF�+�E�����wS�ꑿ��W��_�T�)f=�A����u~��o�:&�%lW>�@W����=�  ����έ��Pڳ(A��q�FbP�}κ�����̛N�}�8C�&ypz{�UQ\�J��x���b�B��΅I)5dG�G�]WS���]7*F9�7t�����?�Z��A~�i�<}�͒�)�J�󌃔�K*iބ���0*c�35e�%oZ��_� �@��s�ｺG����gwr�p��D�B�R�%,�;%P{$w������`���A���A�S�P&�ԭo����1	�����0ru���`�W�d'��#��!|(hO`�šR�A�^���y�q��8�"a�EO
/k�<���ȕ�T&�C-�-c���o�{�{4��K�������g�����3ӳ�BrU��N8�>���Կ~-�Rw�*!�'���P�H#$�8�A�θ�r�y
�����[@|~�i�2�Bc8�=�q����X-�bc��	�/=\L��HSE�Ga��.p�}��Kʈ?z�G�Z��#K�Ϊ.�S:�W%;�|D�I����P68�U�;���0s�a����@Z¼2`�)���crjB��m �9�,���~�����k날�[%���߫�Z�y�Ù:$��p	�ڼ�%����ُ"0p	���?+Ȥf[�P>`kI	k�Z�������pC_[�Ԕ��=�z_/����J�K-
�B�;o��WJv�L���u4����x��'W+=M%�;�B�|���Q╂P{82o<w���ϛqo����.��W�޸��N� `���%��[��yhBhΟ���&��I���le3&=�"Lߚj�>���v����toR>΃�:v!���4<	iB^����O��脤�f�]��c��N�-
Ш.B�^�|��3� m��H��m��[�=΢�J"��֨�u��3C`~�𑁗TEL�7ϐC`O��kg�bi�J�A롃3mz5G�(�DN��؉�x?̘�����&W����D���aH.&׻� �'irѦ=,T�����*N��T,���I�۽�����,� =1D��[�g!�������i��{t�u��e�4�Xp������U򔝵�,F��*�H��7Ќ����	��(Ec�k˕�k�Ugq���t���`�4�靣���u�N~E �R�'���H������q�`j9�g͑Yh���\=[�W��O�"� �vD�4p�X@�q���������܏eXO�Ysc�SXLa�ԫq�2�4<���
˸��F�~��J%������]�����Aah(�'���צ��3X�{	��Y�]7�_ݼ�4U9���)�P�2f��Λ�G�Y�q��o5j~@�H��.��"}�&l�~Y)Ƕ)�0�+�E�2�x:�>��q`�Tu����+RW{��P�t�v�>��e<de�D�=�����m��M{8����ZR���}�� ��`;8�j�hoU������D���V�&�n�9�)��� ��Y�i����퐫���`(��!�5��"�h��U"�P�H\�j6Q�� C!���%���&Z��q��0��W�lry 3v�ML]4-=/�fh;Tn�3�3����ĤB�������ͼ�r*.��-[���a q甖�Bs>t#�(sȜ.��� �bH��;fӫ?�M��Ka��F�֯����7?�p|��
iJ�r��!D��O�(y������o�g�����?��<o�]���t�Y�K�.E��k��+�.�!��t�k�%t��$�b�E�Ay�(���,�W �$���������X1쮹���9��-z�B������t���`�^}Ż��V��2E_�Oi.A�j^ّ���$������ǝ �Ά��������i������͠
��顪?��C�˩��ߘq���q��V�+�jd�2g�����wB�:���Vͧ��vf�2�L�Ӱo(�墱�F'�b�5��?4;y��ޚ�������,�>�9�LGd��j/��z���a���Ѭqy���G+ќ*�0�IGͬ@���p�~�}]afIhH��j��,�j7Y[NBd�����b֔&Z�+�?rz�s$hQùdx����R
AgAW�~�iUlHd&�t� %�}V��-��p�� 2cu�M:���n[����-�X�,Ψ� /�J��ӯg��.d�p�5>�j�8~�_�$�C�mSc����o�˜�s�k`{�e^������������`�ƂG�Uf}*�N&" n�#���&�k�דּ2��s^�c�C�	πK�Xh@HMrM�^�-JUp9Cc���ڵ-�N��Ω�+�=g8�q�p��1kI��<����@�?8FUPߘ�B>�_��Z�
���t`?�rMN�r��0͔�գ�Ac��	_,�(�)��Uk������u�㩗��
]ߒr���M�*�j��@zZ-2#��b3�P�r5��'��@��i��9�sm�E�>�&�1��(ޱ�*y����~�e��l���R�9�s�M'`x�~y<���nNN7kMb0}c���)��.�javI���D�1�c�C�8c��Fl��GܾP�����n�t:��U�,Ϡ&A.��ߠ4� T��w+�st�<`�|�x�{�J��B8��4�
��;3`q
�-�K��b��(�3����H �������Ԑ_���v����h�^�Ξr���NaH�I��>�A��vT�$o�0�} ?k:}ݔ`Jp�A���JOJpx�鍊�*����!�4t9Cy�����G����@U����fj �da�&O�D���6�� ������}GR�,"=w�e�\�	^_����s�GdyϽzn�A�1�c�mF1��ь��heN��5�7���ᮋ�����Gh�x�f�ς��)�<;�E��SwJ�sڴe�+�F�QG���k�nIN	��xj��9k�i�B��b�h��s6�u�u��lz������*N���b��`���#���G4º�5͐�f��������6��~�Ȳ3�)��> -�_u�/Y���$_�$=���6���?���ރ��7�=����X�ޞkQ%�f�C�au�y��WMF�����1�:G�1�O���p}�`���\>o3����D�c4Yy�:	�?t�1m�W@�҈��"����A�$�'�ʡ�p�r<��~�(#���Gr�r"�D�Q};&e�,�E��U����j�'~�R#�`�94&V�@�!w��}Y$����U_��T�}t�?&s�{E�0�ɭ�L$�r��^F��"q�sm.��+(G��L�����5T_I;���#�nx�;*5�ҝ�o^�s-,�2-pyA��=a�>���Z�S���L:��V�S\	�p�_G��Ţay�B�l��6>��\ �߮4'S��Uїṹ5���h)�k�8��۱�!B0舻����Ύ |v#�s�-tfk�<��;b���jȮ�<�Zl�C�Ԍ����S�P���ϖ/l V�l��@|�#Z����o߽C�W9��*�2t_�mzM����[]���?���'*z�*B�i�
��3r���@d�`� \�������dt��`M��(��%�����g�@6�����D�ĵ(�3�
7�rLTIJ��bP�h&�()/Z~�˦+��hZ��Uۮ�b����6`"?�<+>�b����C��̜�A���*�L.��^s��z���g��[�gv��͞i.�z��\2
E�&�o.�z�wy,���Ʋ�.Ўo�	���x����}l��pK�E�pK�ç�@�C%�g��hJݺ�U�2��L��V|T�fж(c&qJ*��#<9����p�B���:���?}���P��k�-s1���Ok9�DwR%���|��ܣ`�pG^�/�����sN�U��"j<�D�:��dV��r7�������EҪ�a��+�zC��5�w��'*Yϲ^꟤\�|�-K��������LLY(M@|�	�B/���e����#�'.XY��fH��2;U1����K�۪�h�
���y�N.���ђ�F3��څ�i݀Ӡdha��cA��.[=���g�L��B�w��cx�%�v�I^��a>Q0��`A�[X[Ң�A=E�,h����S�����M������%� J�`�?���������Uv\�R�6�OV�nH'�2D�T��i����3D�����^ٿ��4�XD����d�Y}n ԫ�U�O��[R�G/8'ʑ�]1���/i��dV��\�yZ�s0�Y��#�+�������C��6�����,��M�X)���Vθ�^�t�YE�l�>�������{�A<s�nwGZ�r)Hy��`t�5��/�i���G�^��J̿��l�@!v�}�l"6���V�w���1�d�2 :�����װ=�'Lxuj���e`n\���^|�<��X�e�s#���k�}�{���c���e�j.�iP��kS�zBK`��)�����5b.v�X�{�lq�H��>�fv�����aja�}�G�,��g
{�O�5���"�I|)��#���W�5D;,�äi�po�2 ��
��js\�fQg0��c<�x�����-p�����	���z�שp	�+�ߝ�,KqЯ��f�����VNI%�F��Y�W��O�W�`.>r�ͻ4�'�kPS��s��,�t�x�I��B^�쟩�v���/pD��˯����<�)��U�D�Fm��xJ�J�0��Ů�li|&�7N�hm��5������N�O�Vo-r�O����nȾI��w�B>� ²��|8g]�.�e���D{����2[Dƞn_�_� �l���`IJ�Ƀ���|]�]�����b*1$��4��+�|�$���&HV��R*���0_݆��)&�������;�K��uRI,�J5��?�?���1�Љ(0��W���o�y�]Р���B�1���翫*�dA|�����
�J��]�t`a־*rv�5��ܟ�3�&E�-o�a�����z.�lcu۠��HL:8�'�nʢߠyR�Թ�x��i,�u����]d�� �c!Q�l��H�2�d1a��Zy���yj%����ǝ:�iO?��[W^OH����%<�s��F�L�f.K�}q�ڨ��T�g�'2�k�;	E��R���g@��*��Y�A��'��@H<	��aH�V<H��f����^ω6*l�.��3��=�a��_��	l�C���NH$O�x�~a�$��&vC��D�1?Uo�Ő��+T��@-Q����6�S~d��\0�ȥw�Cj��JmA��X65���cQ��(n▷�|����g��3>����'6�o�^�u�B�O@#��JCz�����z�*w�TiVL8l�˚�N�#�uF����fJ��Ԛ���.��6�)^ �D"��FRMh$�T"Fg\'�%�1Q\��� �S_q�g�eZn�>��v^V�{V:�,a z�nM��1����ax�$_E����f;�k~��}C�X�ղ6ֻ�Z��$�CS�@.��D7�)0��r�M5��;����[oO!�Xqᭆ�t�-g�b�Lz��~�F��4؄��t�w�f��N�@y�C���	��s�u���-� �ܓ+�0[��[Si�����O����"�.�T�}-��?hʖz�B�����	kh�]OIh'������`_�$�ОMt�8�L�-�1�l�����37�5+]g����AA/�Z�ͽ��(,r H�(�� ��E$�IG�k��%��qAK��&_Ʋ��V3,�d�˛��O�C�&���q����v�$~w���i�e��م&N�ɭBv��k ��&%l���9^�A~f���,ץM�tT�;*>(B����(����A�W�V��T/����:A�X�T=��p����W�����)S^��H¢/�����$�6�$�t�.�ek-�]�n�ۈ*�ó����q�oT��ݙ��Os�B/�ֱ?�a�;8#���8zs��mw� �!�9�
���wR����IQU�_׹T,�y7<h��� ��=�S�X�6��m���{-JSq~�2A~�y�;�$��w�0)L�K�ꛋ~��=9-%F��e�Y#�'En�aS'��C;�~=�ހ���t��ccj��Z�UWX]�<�mY�ӜZ&���������߹c1�L��1;��8M�T���@��Ѹ\,׏�v�7WL�R�A1{q걝��.Vx�m\�_xk��kJDZ�ۅ
�E
lϷ[�i���o��GE�(^���x�������V��O�E�eb�T��Y3�j���/�f<dY�m����@�
���H!@XK*�^y>��s�/|�wj�*�?���?9*�(nUSA��C	�P׌���SI��n��U���M�����Lv�yG�3�nGՉ�P$> թ��{��ԟ��@�+�
��#�_��q_\����:�a��m����A��j�+�����Z�;�N��`�q��O�hu�gc��!��X����9m��F�c���gM��3�Q�jCn���kHR,�����ݔ���K�@N޹�آ/�jo� ���}B�Q��ǋNː��� oi�O��!�	Hų-9���v]P9��.H�r�v��{G'����t�]q����zBNQ��K!�[Oc�bN�5e|�ڑ����8l���2D�+���y���E��
����b����N*0�˂r-�%�����N���ψ��S��z��Nĵ��[��z;�	`ߩ�{� �����3#�O��	�7l�:6qnv7��O�э��Z�=@�@�������_B�M��1$ͽ�h_}$S�.���뱄���1�VK����j���zgУ����h����X��@�@�4璸�.�������)`P�K̥�D#ū�<�5�u�x��X��\�y&��M�r9"%F�q���Y�lFrҖ�|E{��]�w���`�;+�=G6tcz����$bT��ug�3g��o����;֘x	�M��au�����i����{l'E��ɿmZ����*�h��2�KE$�J"P��KF5�^.% J�!&��>���}t���k	A�ZU,<ü��[��3��9&Ԭw6��D>mhVîp���x3~��A�G��j�+
������^�m:E
.j�x��C*N׮>^��w�	��<�h:q1ҳ�	�l��:с%�/e��V��yh����� ��H�=�&X܍���J���IH]�A&��>>v<�N�]c�QK**��Fc���	Z�H�%u�4~"f�I�U8��ԸDM����h�4&`�"�49�r3�Y�ʅ�Y����+����X�(��̖ۘ�����.�V�Ď>�&Cg��1��ʂ�@���90�cZh�I�7u���S���s4m�����2�mE޷�&�6	�.2)G�^�I�������(6���-l�)�j�˸I�(.�� ��qB:T�Bw�vH�����2����~�'@�����k��_�f�[��֖�l�io�j�N��]'���^��`ɴ����V>�gӃE:����]��0ɟ)�����=#��z�o^m�V�K��&��#&���0𔈤+8��	6|�H.Z���хc�*��Uf�(\U��n��~=e��2%�h���u��N� �W>Ω�,O0�I�U����]�t>�o%B[�0�rF}(׏L���OzR�j�[v1U��b����Yl-� ��qi�jhJ���u=
[�=&�n�K��,T;���)�D���^�p
E��'�@�§0St <�!�n!bau/n��! §�fh-�EH��<�Bf�<5���TELib��i�(H�K�ư�����k��W%PRYx~�ݲ�^ ���u>�lT��(ƒ:j�5)����х��'���@�`�*O�Y� ��qI�1(n�҉1�'��T����z�(ĜCͨF�{���k�zZ�K��~�ő5�@B���t!�2é9�i�rg�F��������ذO,�b� ��.5m<�H�d��v縜�[$b�Y�Q:��˽-�>lZ9f��\��]�z���o,�� ����F�yԬY���݄�]tF-����:�~V�GF,���X|\:�:.��Ū�v�/��S�X)Gf��2K�fj��e}S�p/��k�H9�ٵ/o�^��Z��b��b	����ec]dKkmm'��O���SD�`Ҕ�WTo��gC��E1$Ah�]�~�q6�,��Ǌ���� �����Ǡ̵��*�f�����)��C$�[�gT��G�Ҡ�3E������ ǿ���LT��̍,�����-h�(!�95���f��bV�3
/^vC�{Xq�TA�{�06	=ZU���'d���o��W���{��~ì����bW�
�����H�RWֵ�)q�� : ͘o�ѭ�i�	1쉽#.*`�mN�F3�k��6�A�C�H�2�-�"��(������>�9Nn�+� ¹
t5���D4PR�W�(����J���E���DN��}���v�疏<��xуu��Z~Fm�2�Y0�cmiG5|D�`�2����i�'HoWI�	˪��k	�:�]�pe"��[_�ߴ~O��hwT�p�6��3^e$D}cqTsoKjhI�$�hl�kR\笖�=��Ɯ�VK`�0.iv&�yh�t�p�����F���6]v'���O:W��oR�J/���:�!d L;�cY$ 8���⫁=ytn�d��*�����e*�mE�b�~�YL+(*������]��	����%(_*ǐm]����t��>ޱPoQ@�����'�#P�`��Lƿf{���mxy��&��w��cĀR��jP.�Z��YT)��W�ż͹���ʫb�3��GZ }Q��`)��k;���$<˝��mi�:ҟ9�_��6���jU/��W��:��SƄ8u��uq%�8����<L���3�X�K7f��]��$�4��ӦT;`�;��ϭ�=e��A&�d���R�3["�Ir�������dy��f�n/���:������q�5Y�"~xҗ\y�J���������\�m���M-���v�@	�e9�l/!( \�3��N7Gi����ܬ`�i��������4#)"��@���nYg ;���*���u$1�S^�� ߭l��-B�sWo�fM�?�W�d���^:SD��O� ��u���8�3^�J?��n�a9X�����-c|��L0��(�г]��KG�^��Yd�ފ��5���젝�_a'a�]������
���g��R�ݪ�jSZ�o��N�����>�J�N�]�v%����]d<U�u22s?c�R��ג��pC�n�v��8�Q���ݙ��.נ�kN��fn���M�9�����b/\msǌ�?��z��CeO�-Mʶ��^5H0���NsfHa��rm�s�]7�n��\�\nzd�VԺQM�u�P[_Ɩ�~�yK��d̋�)�ۆwWNv;��t�<�Q�w��3%K�l��`�b�.�!��Qmz��3�_�Я���׻�.T���N֩X��������@�z�����9�ӡ��u��l<�ab4���$҉�:��b����*���_NO���f�b��#�X��17/�4�փ�w�C�c�&P����_RɉZ��uitD���_}�#�m�=����JD�nId�W(e�r�PNA�<��N�-X�a��\w�����\;(ݪ=Ή#C��f1�
U]h�5#<�~a�G�Tb�w�?=J��00�o���W��.���+W0�Ċ
�1b[����.L�Ju�P	�6w�%���$C�&�[/!�̱CC״Օ.�$���Ir�����Q�b(:E��=��Od���8�\u�t)�z�&m������j��s���H��S��c��K�K�������5��"����5�=a\����r��`H�1�6���	�g-�"��>��7��2���/��r�!}�H��#��Q� ��7�����)'[�=�^^�,>O�!��a�F�ʪ:�0�y���]nV��k�\�?��sS�d�t�DF$�gRd<(+���m�gUP����'a�W+6��_�>q�� ��H�9�XLB�Y�����;U�j@�e��d�[��H(������W�s�Ճ!8h�c�-M��k�\�ę���<�e��5x��ye,u�oOZl1���oL@�`o;n7	c��{��e�k�Ҏ0��+�����W!4�����O,Dd�4�@�0|����6,L%/&f1��C(:�N��D	C_��ef�n����s������ �;o�=G�d��$����K2IX��.eT1n��b�n���lׁ��榒D�tJ�J�Ly$���i4���w*�w�B ´)kS���b]��ZI�! ��M[F}��q��N�4�a������ڸH)K�{0�ޓ�	����at�Lt�7��x�Ӏ���7+� �Ӹ�4rW!Ǝ��b�)��q�GD�G��M+D�3i[xe�l
H���=��i'��`��ί�E�-R)��6�Bn��Cʌ��<uy/�{#.r����߅o�_���ʝ�s�����o����j��c.j˕~(�;b�I��Z.��crD�8�lӊ�"I��Cq��]FT�>MX�NoT� l��.��Xo>�(��=}��� )�G���d7�;!��jm��L�n7������+�եo`��h1TY�� �����Ǖ�h�P#h#�$--��Z�_��z���CEL|��?4�nѺ�2C�"􎑶�b%�]�#^zmP���.�B�����C�����)��ȋ+�Jp
�}�o�@��CƮ��܍=7����4�I~���=�^�u�{F1~��Jb\@f����0�R�C���/!X-i�곸E�h�`�W�U��R;I��(qk@
ى'�M(��!0B'҅|�qܔ���7���H��P�:��J.:�_�9U��o��%ǐz�Ṫ�v�5���N�Bh�� ����"}�������Vs�㊸
O���L|��3�f��I�b��h�]�,�.'��|⡚�-g��(�NM���;�_4�AJ�4��/a�3�&>�w6��i���r#ӌ^���>ߤ֓B�Eﳐ8�� �@{�G<d� �_�/��a�Z����Le��C���O�^�V�Ua7��`�,�������#w��c�v��� d��6�����B���&���M6xa	3"V0�~��Ao��e/4ꊪ�g{qֆa
��)4��"��n7�m�~u#ى�_���{��iS��ɴG�I.����(˚:�h
4߰nw��ϻBJ�w��/eʜ+&z+��3C�������hu���+7ĄPiGIN�����
X�Q�31-7�3U�75��5���uoK��%�0C�'�]�	}9bO��Q"�r�g3.c`0�ڱQ����;�no���, �ľ��������������zf��������*�� Nc��~AҿzJ�L�M�y����DY3����
A3�kpq�ϠnG�|��C}�-��,%b��${�p��:��+�'"~ù�d�1%&A*�O/�`![�p� ������ǡ��4�d�A!x�kԨ#��@ʙG�zy�D�K���%�[C>��K�*�G ����@�u��G�>e��.f�틶ZS�������,)1�� g1�?����Y��5"�2�ve.�2V��݌���y�8�W;�x���Ϯ�o���]F*���hN�RP���� b���_˵�I�u�/ɭ|��2�C�����{�uXxHO~���ox��oNV�]Z�sY�`Y�݃kȺ�IEχ���.$��u�e�T4�k���F3lI�%�\ FeE�6d��M���_d���I6�,����=�$��7<��4~g��Nc��=�L�ؑ����{��/ ً m|Η��|�>-��@�(ED6�4t�)�A�������F �ג?�-���ิ����O�_M�qY0���2�t,=8Dby�ӘL��)�,�,�ǀ	V��YB��$��Ϙ�����øO60� Á���#����h����K��d��Öd�@I�u���{�G�<� ��K��>O�:	�Yv�+K�*&2x�e/�O��1\/�,Pp�3����~ ��r��y�=`�e�8n2k��4�3V>8"N����A1��h�lOQ�ʔ9��M�LǇ� ��M�L#S��]��y����w$wd�s���0V;�m���w�:���
0�u�W:�A�ÖxqPص�%�ӫ�fH���@y���>ݏ����θ�9��Ɂ3��jKܟ�˲.��	�p�d�a)�>Q�x��%�1,)���(d�!�e��nŜh��\����0�B��I�=�zx ������$i-{-�ܬz#I	r�R>{����p�Tk��{�v]5�}Ȧ\׳�0�����rq=��WR�1��X��Q���*}����*q�P��˓�D�U2���/ei�y�m�t�	!xF��K�sy߲��`i�n�O��G�n�816 Rc$'(9ed����2��t����� �BS_�GS�8@_��/�A�Kj�4Ia+���r6tu�s2	�v���L7�d��PC�����ݥ��0�����L�{ui���O~1"h!�9n��a�}dmv��4^J~'��lq��s{,�Q��ƒ�0K[�M�&�a|�?P����:���<R�������®h���ؒ�Ŋz���n0�O��b�� �I�7�U�3�epj�J6"r: ua��a���iK3�߯>o��4����-�%8[��(��=�L�59�����d�;���6�;��i���n�T�%��
�4����J�GePI+6��k�]��8N�˻�m�W��)K:k*��cP!-����^?���A!��>�U1�7��~ͨ�����H�K�T���ѥ��ƾ0�5��ZF�S�H �P�-v�{�G�n0��t�M�nt���g�*9������'�ɨ�oP\�.��+��n��i���C(mB1RZ`4Dp��EE�[��Y��^��I�A��j����a��5��c쏽R�q�	�a44��	ZF��)�x�8b�{nteyc�=�+k�8��
R�:M��Kl�mqs7�J��Ij^�D��V��ѩ�+��鄻Bíh���5B���r+��=^�s�xem�2�o=(Q!<Y�F�������)�4��.��[M#hW������p0�j�V�:a����k�)�����OFm�����!.�RNr����@��@���]�d��:���u]�%��(C��&3��D����!�RA�z$8bm��,k�0,l��c�ie����$ ��i���XM�Z��k�(6���t"~<���y�?��Q�	�D�{�M�[ـ�#k��J^Cs����q	[�%;fc��%��%
��)<M ����Z6:~�*��j$��ϸ�j�ɛXq� /���G�9��77���xo�`f��� ��7�婃�����3�c����t��Ԣ)#1;/��P���s�ՈB�!.���Ex->�{�ۚCZ^Y�X�>�؜�S����3*b��٢����6�,�})�g�X��'����SR���3��(�'f�JI��7�m�}���Ah�͡E
�����͜�7��
%�/�]Bp�$t�� =w�΢ 
�fU.�)�.b)%�����P'��)���R�=�YJN]��LK&M!ߒ*�)�U�}��\`�Pؘ���إ�&�s�=xia���$����2 cn�W`CmzV%�%���
��t�-�Q'V��T��H~�~̪� ��mG�O�Y���a�)_��c2�!�<0g�m�ze� �h8���(wV���퐻|x�G��H�#ђ��{U�ǦB��׀�"��kӮ�٘���F���<�1� bΗ�̄"��O���(p�l�q3��ȝTP�� ƿV9#���~jݪ�v�.)ffa���#�ӕ�u�o��J��ںr�Eޜ��N~[���4U���}zZ���ZU�G/��׬\lrrw"o�C���[a���X�87'cs����-�Ђ��D�F��E!�����,)���8q���D;�{IS[�䩼��J��'ҟ*�KK�KE\:���'�Sd��r�2
�
��/�)+�����/�����<3v�~{�?�)���;G�c����d�)6k~���!���
&�=ab���������'���#��S@e8c�[d�])hT�Hel��>As]���[�H���LrZ<k�C�rP���I�1�6C(�S�Z��^"�/�)/�w\X��o!�fK~*����\�d��3)v�z(�Ü~�l����L���TE��������{}z�	�)�|cvH�<��;�ja��[��Sf9�EJ��8�x�~X���hNL5l�@�kv ��Ċz�?*b;'� ����汉��}Pͱ����ط�֚qjA��Ɋ.��5���c���B����CqC~-���w��įd�y��K1�T��h�۬�|���*�sQI�u����:u6���'w����C��c1wa%:����C�(�TJ(ܑmw�#q���Ee�5��(2��e��+<A�9�+j�����Ȅ�R�/I���b����W�*h]�l�K �r��
�v���^�4��>@GY�:�#OsR�F3�B�����m�Y ��>&�X�$�t)�z1�0P�_��z%�@�Eǿ�r:�?&�����WtUl+9���1����2��lm���u�V�,�OWh޼���X�4����9a���蒪I�X��5ь���*$pQ�uC���a!� h���:Ԇ��4r�-��ɢ��rah����Q>�*�	��\��X[p�����Uk���%ԉ-�+�[ �����]���P�'�%�F|w�{���s�� _W�/�s2�$�<,�2,��Q��� }M���wyz��+����O���(�G�Y�v��>ҥ\��b�3d�mH�bŸ�(���{�ajӸ�8R�ThD�T�[�~\����̀om�uQ�u�h��]���DT�+�| 9�9fwL�K.��J�Μ�v��i�)���	V�,@����hu.;A��M�A����� ��} �j�K�ȭ�A�)�A2�389~��b�@�U����m5c��#0&��D�מ��.?��o^�,�$����N&��O�G��Mt�������t��3�}�b�"a��G=w��CF��ܼQ��h9�)���$\I��z��%&��ؒ�4��2d��6��*ی+.��p~��������b+�c�tL�RT0W���/�To�q'�g��@��~�I�us�/�_�$yj6�c1�I���ճ<3���n�HR�8\�h��@&s-U��[��ԅ��R���	Bͷ����ȋR��Uq�#��pG^a2�Oa�qX��hK
�oˬJWO�@�z�f�l�ŵ+I��[��#hG��X��w#Д�Ɖ�T&��I�3E�qN�e,�a��B��
�x�g��� Tc�?�e�ٕ<�U�p�����޽������ì�͎��3�9je�02]B胲��r��Jy�yP�vo=^h�e_5Y4�*,��j�M�����Mt�5T�g{$ʍ�r�6L&�"*�Ɉ��� �ۅ����e��
�L�aj���B�i>YI���v�6p�ޔ(��������w�O|~ԙ����n�b7��h�u�����n�� �˽ ��LڬO5�5}È��Z��,����YH�Ou5���R��7&B;�E����k[.*��������&:�ޭ�05���\�Y~�(���/�^���Q��Y�M���!�������p���E���p�˽/O�	�Y3pٽ6$jWGE�e�A<�Q��A[�ʵ�PS!��M`���i=$�Z­x�T��T��[oB��u��Zq;
3�d+֡��&;��\1�Z��q�����'�T����cԨ4 �cd\��t��uȝ�b��͔^����i�r�i�ء������1l�/�	�8�<|���G��(q�Q<�f��yXז|3���1�2����~��r�gso|0D��^�i4�V��-k��c�J����v �ۤ,�\�}1�H���{o�OJ�&������wl��NKQ�L�� �#�Ѳ�HD	�x����-�D�쿖 !#�t�ό��#��w��a��B�>UX��.�J�<oݛ�hXt0jq�i7���}�D���,�0�a)^?�*~ө�3�z�`m�L�'���Л��A+u%���*�sK� ��g����㓺͋�N�?}����,�q�F�ws�+N��Qct�dsG�"�$�\7#;V��p*�![��0������#U�?d��l�Ԛ�cT��c�?O�GJ����z��F�Ǧ��VC�tt[)���a횴ǥ(�K�f<V��$���*Nd���0�r�u��Ou�y�؀_x�nwv�dK%�p@�Z���gh|ݿ���q� n��y�z�
P��#C@��t$|D��ŏ�;a?��D���$F7�h�+w�+�o�������Hb[�E�گ6�0| �wqo��,���\L���1��~n��t��)�@�����)�
G
j/��^��Q�ghj�^+-I�&5�~�IO�iPYS�ela���RW j��wN�8*%y�2FI�����u�ͺ�"��=��z���b��w��Z
�rj�,��lyeA�����F�S$f˽ކ(i��Wb�,�7��F���\>�FY�\���-����y�@T�tP,F��Y���x\%���������sng��~E(R%����˩�0.v���[K�"�Y#˱�@�M$��lA7��Y7͸�⪟�������滥�4�)�o۬���}Y��(t��,С��z�
�ק�Ҽ[�T��͢˧���~����l=G�CI��&�� B�Ә{/��&�/qB�����-�����%��t�I�LjH�漦͏y��^�%OZZL�0��{f�Ͻ��X�<Ő<��a�V�4zZ�<II<�� ������D/>���5u���}p�ͣ������qWZ�Q#8p	z�՚�!�qkjS���A�r���u(Tʶ�Έ��70�����w�_S�*�6�KW����:�ȉ��郋�{���h���N���J$��M�Eܰ���o)J+f��3P3�_�'��6��^M�}z�Ш���`(��ɼH�
���1ȵ.��=/�Gw�+�����1i��B��JA���5G,*�2����u�N�\ ��@c����$�b�T8D�ڹы�"�� ��t@���t�a=��S�q����f\�p��&�z.�R��erC��G
)ɆQj�ڭ�Ճ�mC߼���^g��>�!�zꌴ0Ե7$��2s�����u������ �0�`�7�G�հ�髚�x޺�������� .4��Y�����g�x��pѕ��}�:T7'�]i�|��z� �϶�+�{0�Y���o���(����������|f2�zL�xWɝ���ֿ�`��n�������x�w807��)����z�lM7:�FI�>�NL��^=Z�}rA����>R�Lo��?M3�5`�ҽ�MAk��k���I��YE+����>��Ć����@>g���)�ZG_�^��XE[1�.:uGy'�	�LM�5�� �3*�O���d�H��vT?��h��i� p�#���@�����Ȩ }1�c%ۖ_���8x�y�ҚJ�5�"�:��a����r(��A� ���^������������`��A��Ҏ��]����6���oA�U%���v;��I/`x��b\�{톐�m1h�I�
�/
HW���\�CA�i.���޷��fLZ�k	T)��&xM�S��#~4�����w枭��=�C�8/����Vy`@���Rc&g�q�.�5�e���[�p�bo�y��@6�qvk��8�l}pF@S�'%��(=]��&�����C�鄣%��!�$���N��չ����u�j
�����=���|R�O�f�K���ԈBP%�`�E3[P&��MG*�i��7�ղ��_~K��U�;��ɼ";�}��Fq]��1���O�*�6��c89G�A�s-q�z���3�L�5%��AV�v���i����R���f�n����}D9�F�y�ON�k���H�l�����ئ� "�$47�(�&�D ��o#C�����>�r�`�u��1��X�<T{���$b�+˧��#�<��5]Gc&r����r��hY�uQE���g75�Ji����%�zհ�~p�M������x̒��ve���u����lO�z�e�KA!C��IA����~�a��7S��8z:1�Q��7!���!m�?p��!��#�e7�8S	xh*���d����� � ;;��� ����A$z�xdȷ��n��ɻQT>l *�s�kQh4r��^	�3��������wdO��+��������-��JW$���A$�(Z�oF"�2�W�K�zEEB.c���P/��١;B�^����ŧ,�܂��4�ƅ����ȶ}�c�	�!��O�D�Q�22��a���-3��C
8������Z�gA�?�fz>��_���x����!���·���9���s��G� ��s�LT4M{d�98W�Ս���v��v��"g�(Ϧ�l=�!�UeC�����A�p�l��Ly��xxA���\<���ߠ���cC��n{�Br������%�;t`IM{�7���:5��&�����J	�z��-tn���Q������r������qn�c���&�NM�縘k;Eu5�䢃����#�8����*�հ�{FzI�n�a%�g;c�ğ yǢ�\�L��0wq�.�9}�����@��RP��X�?_��#��.�nr�r����"���q{1�8M�|ʴt$»I���'��+e��wG��� �3���l�9�w�+ݷa6�jNQ�`���r���F@C�>�lbk����O V7���k�ꗠ���&)#�Ptn��|	��3G�u�x��!����S�;2y�b{��0{���$�hS�N��������׺"f\K3<%x���36�;k^�UK�����`��K񜁛���u�&��Y���Y'��ea��ڼ��}�����	&'MaG�@~j~} ����	p��C��b�a����l%�0�G���Њ��	]'v�q!�g@#%��5>��Z���k�x�R�N b0��`�G&uAg`V�8U.f��1a<"w����aW
�X<n���
�*�rOu}0�?�|XS�Z�a�^��3���Pj�!]A`S���gH)d��DY3Ea����2�=I$	�\���t�;�����V���^Ɣ�hv���@�q�ݬMU���+9S�5�72�}?��A>�!��Z�]��Bk���^EU�qG�s�N�ۡrC����+�y\� b��G�)�1Z@��+=f�v]iג�sY�=�u�Yn�h���C�:]� �A�\��/�4 ��̒��
Zt��-Q���MdN�ZX�&�K�p&[�V���<��+�d�����"�&�/���/�d���먠&VzI��l���Z�0��T9��[ҥ���u`��K�����-I	򍬦ɷ��v�X�TR�������L�'��n/%����U9{��y��/,��.�S,~z��#� ����3�Y-���Jv��c���LT�v�ZEFN$�h�}zem�G{�zd5DB�	�;���&u���x6�G��'s�����>�������-��_���r���
�9���W�n�ՔX�{4�oVo�@"�7�mJD�7�cJ���Ľ�E��B��T���R��C�N.A'��PMU��}rtv-�e���L?Q��Eί�_0��y(��qk�	��KcY�'V�:�N��ug��kG�17r��he��4�u�5���xv����~�6\ۘ���h.�z{�:���m�����f9�������|#�����*9����Q���
.p)o`h�$�t�_�H�(�Xh�<����f$��x�_
���qF�̒f��./�<�o�GR�r���Qi�܅�}���_��ƻ�j�\@ȟm���"Pk������L:��B�C��d'��!Y��g��	x���*�G7�1=�2� P5"	����Jv�E�I���j�+���Ȉ����;^K�O�o��gz�� ���o��_sM>�(�iEKJ��ދv\󀒱��Y'zt�7�����4�}��%��3�N`�(U��;QHz%}�h�T+O �&g=���S���L'zA������}z�(�#rĜ�G��}a���o���0��u�]���vzۼa�#��z ��DhlЅ1���Z_�o8@֋�'�W{�t\Y�/�5�	���mEJ �^�Y�Fy
0�Щ���Ĉ�T�&kR�� �nBG�� G3��KN[?���`T嵌�L����{"��㲠��{�
��#ZO$����?�,@��� �)����H|���x>�o�ݱ%)�_����	^T��2��U���م �o�xb�g�'UB�6��㝚�~�ɑ��P���p|�5������y���.v��NK�����0���3��{+�e��.<�w�b?�O}ᶊ�uq-���mr5�"�Ica�T� +W	d+9��g@�  1]JԻ�:�gJ����cI��н�������5Y�Jn�$K��U.���χ�jZ���K<<����]*�zKҺ%��N��	@N��V\�ď���82}����/L�H�=�Y�^�7R���"d_��
��)�{Ʒ��������M_sN=ݍ���1��.��}+wj�58�JiM
Z��v�.ȍ`�&@�yi�\���gus�o���,�=HQ���ܦ�_��`�.�j���
�h�^!Y�+�Vq5
��B��˪����P�l��/.%5H��
�������}�5DOJ-SA��m�E'9���O߼�xo�i�0 ���Z�g.���[���BC~��9E%�ibF��33��~�3w�❄��)s;��Ӡ�����s�x*�E_ģ2��/���F 8h�]���E����ƠΈ.�Vo0-��Fk����=�j�_RMc����!fAwͥ��>e]�ϻr���v�$O�p �w�NQĩ'_�B�Oo�~I�qI�x��q�q�x�[��ٚ�h���f5��Q`�[?{V�!��!�����p,r���8>�m��g{ҵ�&��#��]�vU���LP��L�j~��{�>�1&dǦ���I��pC":���1�#=�)l�2�x]a���見��4g���q-m��A,.�G�̽�ٽ��b�k	�j�z���-a�*�4;�7q�:{��ˡV���܉��/�|e��xB*��f�~(�9�*2(g'�����"�>��p�>z�=�M^̝���q2YuV�,p����`�>!�d�P�.��,�N&��a��G��[F��->�"��Y�ye=T_�;펬~i���ȆbX~�(bo. �EX��2�T��aͿ)�p�T!���;�q�7��f�Tױ�pn!�n{���?���V�_��ᨻ�46_Du�+>�|eɟ��8������� =ş�A�9�7�\L`�����f��}��D�Z�H-]
��Mm�qCR�@�i���k��Å~&�0=�?\�k��Ù�E^t�O��o�gPC0lΡ�l <鮞V��Em��?�?M���P�T���K+,����/+�Hp�<�	��%�ga>���d5B�j�����UѫB=4�pj5���\y��V��SRcpY��LQ9m{��g����J� N_��όj>f}����f>�����?�(�e�ӝ��`g׊>Ϊ��`�~B�5��F��WM���SU$��L�Q�q�4v���#rA2m{����Ĵo�҂�zRZ(��g����S+�����-9��m�t��ӔL~^M=�"g&�P�'`��t����2� R��&�յSN�u㇊Gh�A�Dɲ���Q���x���V�-�`:#ֈGC��_��F����x��n$3�Ə���X�E�\Ƨu�Q�̅5���+�׳4�6�Q�s�-�.%�\��5lE�eM��!�QJjn�cc�t���m��u`S{c5���Z��Jf7�-Oz��i�uі�p!:)�qm���m�/�T�/�vy�)^�\����s��I�tޘ��>��G�ϣ�b�/(����	S5�(Y<+�Yv;�偶�o֦}I�r�Ѧ2��E���@�Σ�(�ˣ7�4E*��<Մ���}�Xc��T��2W���9��j6L�s��2W4f��^�hܺ��a���b�̈́;eu�me=��o���._ٺTw�O��j�0T8����ž+v�t
cr�^��zZ��[Ǩ\���/�H�
:���|%��φ�`�<��!�d7߯�{W�+���>\��9����t� �:o���eY���1����ۗ��\?d�d�X<5�*˾�ܿ�(B*:Y�iy2��.�8�B~��,o�m���k-0���Y�� !�{g��&��`fٓaT��	�z�\��J׽m�QBD��p#���1%*�U��5��~U���h}R��+��M*�'� ���B��/�Nx�_zR�^���m�g#�y�u�z�l�j�7�x.(�m��Q�(Ͼ�Bޖ��B�z�#���&�����X��۞σ&��ECz��R���.�1tct��뛃�p.��Y��7����3��K�����?+mV�N�PLc�h��z�gu:R����1w'{!6<��>y�kf5����4І�1�r�U�~�A����]�I���*�������������b��I>����4��,Y=Pq�kf��X9]?�n����WQ��,�Iu�a(Uˊ���.l�`ԗ���汞~f�cЙ�1���+�/ 'X p�3���DM����SӦ�)��Sm��h�����k:+.oε����}hj�l��$���_��2ɣg/qt�=�C�����'"u�ŧ�B���9��\��R��k��F�i�A���� �o'b��� .p�
*��0�s40/��Yx���߾2�r�.E�F��g%Ɠl�鷢��_D�HL�u�;�,J��?���v)U��'�~T���&%���F�	��o�0�dD���B��A�� ��������O�VB\�m��;�����Q��M3:� T����ǩ�:�3){~46��Z"�8��;Zz�ʗxAQV�Kk�&�� �gK��_�ET0�mR 
Z����D �S5�I�c�x�}z��c��q��Ff]	�E��Ao{_�M}��t�����@�������t��|�1��'&bŁmvZ����NdH.�������F?�fU/��[Υ>��A:wُ��Ke��7�]�J���)����g��mʴݯ���ӌ�i8'7~�;�1���uE�S�r�:���yH.ڄIF�n�k��]O��s��	q�7�����Dp��)y<u�r�5���9m � ��\[�~j�(���! �h�`Q%EkA@$�U�(���#��3l,mUB2n~	��Y%�WB�AA#@t�[BJ��>RHw�$��E*��e�.�8��w�"���so�)Yb��딏�p�������!��7�(��hwЃMa���!���w��kX~��Z����i�/q4m\�Sz%��Ch�Z3-0����-���Y��s��_!�at���S�YjJ��=��V���@E!(�Ģ%��l�+�vK"�Kk�|M�N�+��:R0���WX�{��������N��y��O\�A����Բ�'��49`�8#fL3�w������v�긋/K�Kz���a�4�`����X�#�0��L����������pt����]�,�-;m�wTzJ��e5�<j@~W���v�%:����#�k��G�� Wd�]��^�>�� _[������HkyL���W���/�S�(���<�cӊ��L�ve��X���~���'voBnb�S�^'�y����7BjR�J�SQ#�� �~�0,=�,��#߶`M�I���O�Ճ�3�d:�:�!�k�T�2k��"�}��9��P��˦ol�hꮘ˞��6��e�G����uӘ����0f�A�ۻ��b�ŗ��ϔp�w�߄,�����=K{
&���� �I����z�f2T�>�$#��z	 e��QHU�; ,~S%R��á5w�W)XHo��ɚ��܋ˣ%/������iկ�!��С����� ��蒱����ֱ@%�
�4x%;:}>a� +s�+ܯ�-���u��U�a��sL�Ҡ)6���Vs8S�Q�|�d7)�#��F�l���B���\��EF�\WsP����8�}G̛"!��!�7�����L��W���҄ϑc�G�Tb��G:1�*\/���)8ƑM���ć��={�d�x��� �Pg��|��# �W91d&r��[�U�	���L������w���8��i���{�S������4��`Kb�/gO�[��=l�#8�b���:$����7L)�8��C�lNM�o�iυ�KQ�_���s�U��a<�Ǐ5Z���4���/^�)�}mB�W{�I3d��۸]��a�|���R]��)�	3�����0����Dj�P3k�L$�|��Ӹ^J�]e`X4�w��"�i(qf�Ǣ�W�G��T2�ܰ���J�}���p{6ͦ���^�)M�br{�J�],�{�L����IyU.�op�����9(Z:2����ky��u��e0�/�lǇҖ�4vi.̤�݌y�$�.� K�9��1�nK�3������M�߉\��#"z��*�DO���� �F�;xK��:��vv�7�t�H�$d�~�˝W:N�/͹J�V��%*Ly4�#� b��7i�m�P
s�f�i}�́���%.�{΁�V���J�r#���`��3�����+�\����{��Q��]�O/�.A�~�ګ���(�ゅSj0o��fN�d���;�'�SF�V�v�n<��k��C<(߯w&C�Qdwf*:a�}x嗓���`{�:�{�$a�0�(ԒmF�NGxh��:����F+I����4�2�)��C:3ϰDrt `���횤| �m��"��3�m�{~&u^X��w�DXȻH-�e�A��� Ë��4|��85��ĵao �a��;�_
�,������8����M���x��1�ɟ�oY���
N�&O��N�Y�3h7�3��Ѻ���ȟ�&�э�.Mm y�p�w:y�5�϶���<�Ѿ���Ʈ�ȃx��U
F��us
��
� +���jO�UI��Y�`�\��uy�+��%'�pq�ؐ�!��O���H���)[r��X���S��bXM
+ۥ�o�s�>|x�-�ʪ9�Yx��k���i>�F��Y���i@��P�tU0����Kgo�ja�`s,񕲃�%Kfi������t_����>U�,L�Z�)ym�U��#��yz!JL����/6�F3�0|�c�'���.�����yNX�{e(��+����J�6®�<��^�}$�����w>G��IDW���콦��9[ϵ�r�qD���8������Hx������Y�anf����n'��3a&�8�F�I
}��)S.}[�X[�=���k�k��&1V����VL���돕�*m�&9S������gK%��r�
	���ҷ&�N��@��A�����p~N�bHv���|%2:���]Q��%8O�*�C�K+e��O#0��9t�
>�pu8�^%�Ӄ�^��4 5TG�ܠ<�{�'Z�ý���2C=jo���M*�6p �-h4/�f������|����:hSL�J�9_�	����q���,@`����&4{i��� ��i^���B<��m�����^�@�����}{P=�`�
��{���t-8��A�rO�N�r\�s,���t�xp����aԕ|E`�7�`M�Lţ�Ҏ8fo��<�('p�F����, �<�W�w�N��M}�3��9Bn�+3���N,wׇ�`kw!đ�D�V�Ҷ^��'�jiN~ֿS��O#���*���>��~؇bO
��T|��D��%,�i6nW��ro�p�zN�Pb��q�}�PIE����F�}!��wҠXHcbX}�Y��^��:\���{7�K�;&�֞�CcI�~a����s M�~�������g�{3H�U��u�lRR�)R�J ��:b��yA�SwTJ����X� ��}�~5�13���l�C�@�y@7��^w8L9��]�(��]�jM��f%&�:w��O�`u�w�&�z�*���-7v���eR�zˮ�����&��$�\�,ŗ�u|H�_?2~Gn���[֤̕�ӳ	���C�@>	�Ƈ���}���ݫ.�n"/�B~���m�����;��5�||e�^��Q�Ջ��m��2���#��z^�+Ӌ㤹rqM`R��'�M)����Nް�>�]!f]Z��0��/JӁ6u����y^r��v��m�vg���H ����r_���_�d]����Pw���<7h�Eoz;���[f�7GyfH�j�9X�+1��p1ِ2r5Mž�ñr���M�sJ�	�ɘ�Y!��� k�X5z	�k���Nb�~l],��1Pf�dZ+^��_$0�Ы~J.t#�& R����fF�bIa���By�^��,���i\�?��;|8U���o��Ĕ����vf��K�>Q,4����ɍj�{Y����8�Ί�z�ҙ�������&��'�P��;Đ^�X��٫��W�Tߗ��r�l����܃�.�L?
r��j6+3� v
6G��2�� !����p^�𶌋�T� +��}qϪK��ΐ�,-���| ���Ys0gFt�3^��A�ԟx�$L
J��#��bK�'J�cXn�k��%�
3>Vr�V:�HwYS���
VAa؊9W�Y~��J�:{����R�#y!��A�֢�������j�0%��Ө	d㽮n}V��W��V��(��4�."�7�&۸b�vOv��3L�F��Tn3͎g�L����P�8d�m����J���ч^�%� �V��N��2����ƈ��.v�E�f�O����u��M��-e�9�ؒFxW2	������%q8�㌁��gn��ysrb����V�'�q�������Q��.i�B亇&4�0$�)�����hi���Yѻ�ɬ��hߣ7��l��9 Ԝf �����)8�L��gڣE5m��3X�,��_=���<�|�~�[�&���(�{
`ִ�$�[�5�:�?�"�8��L�-'��l��K#8(԰�jPO��t�,V�a��F^�mp���e�3T�Z��g0q��=>C�K���A;�!�ʕ]���k���􌇕��A�A��<�5a�}�y����][�	�y4C����~8֣ٙ��"o���?��5�*�X=�'X�����9v5�����3���7='iUwG)�&��FWwe۩ ����r�e�V�.l�ߤ�jx�*���gsьm�%v�ŕ��x����aA�|�U�|6=����$��= I=�K^t��,Y(.E*x��[T�7�;��{��F����J��o�R��!Dq)8��y;���	���UA�k��~n��~�ޥ*����������ϙ\�J*���5a�/A�Ѐ�c��B��:�▖q.�>IŬ|�;_P�9���կԻ�����h'�<0��5c���l�&����`�5���q�*s�R�@��������d��=��������|���R�*c�g�<6���3�O#��c��	Y�o�aP���W��dtG҇�i��ih �����`:A]�^DW$_�b��7�K��q�v�}A�k��_�:CZ҄�t��@F'���k�c�sRWB��p�|����9�t� U<��Ĵ[Jw��8�m�	�z�*�ckC�mMm���_��N��ci"��3�OcK�=�W��ގ�Mv�O&3�/,�⪢r���ƚ]�z[S����܈J��?������O^\�{�MF���� d�+��N��G�+^�h�^,+��,�����3!Z�<�?L?D2h�=-@($2ϖћ���� ńۈ���C9��Q"<!�v��f�	�z�q�L�c�w�s��{x,�k�A�ژ��k|>�U &��R>=��B(s<BN�b�GX�\�'� ����w۴`�L��t�dM�
�E��F�3Ka���.�i����n�IM=)_ˊJ�>0����qF@�} MκQ��H�\�<��g`R?e?W�8�4����
�� L�77�D�ǣ�IWië���d7�B�f<��H����+~��|6>]Z3��_�w��v��>l�A���S�b�AQfb"oHᥰ �Qd�S���z��n���O�Hђ��Sk&`�EkŜoP�����ުӗKϨmH���J��atcˀ�b2����c�IN��O�[�vx���-�FE�?��z5��;M�Y�R��GU)^�?��f����O+��\۴¼�qI���CQm`�Ԛ��?��ġ�-��n
Lk8#�:�T�p�?��Q`><�[��I�5��.��8�[[� bϠ��.��k|S)ք��(>)Ǹ�U�����z�%cr,şۖ��ZD|��xW\��	|�m��o��ؑQ�)��9�.v�97�KV�g2� ��'1gT�K�r}�K�APB,�3�:�2E�)�Eӵ犷��?�XEs�F�ˤ���ޜ�(j�� ��{����O�#q�wz�����/�F�k%�X�$f��v�����$�����<��u&�-���[D�˕�E ���$O�{�����G�jN�@�ޘ'קN���cuI�e��X�mR�vWd�/�l;WQ<% �q�ze�2�����Ӕ�ٿ���۽>x�0b�ҥ�U��Ü�D?H�O�M7��K�*�M���k����WN�%U��b�4����t�3��y�S��V����T�4�J0]�D-�CFB������ޑ��.�n�����m����y{�7ɖ�6���s�!��_*�Cx�j>�!šI�f�l�:�qޱ���Gq9�>S�҉���ͷ��h�gu�"�BK�<c����6�c�!�]tF�G'WUc������.��.Q��Q�&���Q�!֣V����8��,C�5Yg��:rP��q8K܈P}V�׊M�.;tӰ*��S��3`\.���Ѵ�Bㄌ���/ғ����*Ͼ�حxl�?���艾#��Ϯ`�V R�+��i[It��L�Ӹ:�Z�(�b*�_ <>6D�8+�s�=r[8���g/�gbh)�.�҄$�<�g��]��t����9���|ӆes0�v`�3�辱�`� cɪ��ɥN��^���J�@�̫�K�:���f�C���~}=�v�a����@$��|U�i̔������
�ES��{�	=��7���E�0yp?����E�u9���[	�?f�С��ܿ��� /��s�MD4;�Wk�� ���'<_��ӥWCj(l2ST�9��E����� s�A�0m1�'��u�:��a��'?1�L�ˈ�c�=һZ������+3��x#�b��p��2uh���"�-��#�no�D�v�5;V�MN�X2�j|e3�^gK��d����Wֲ���<�����b�{�$�
j�q����j9�϶��o�| k�5+2C�\�� �#j(R1FT��~o� ��M�Z�ȗ��!*�����P�0]gHPk;�ұ<�[wt�Gc9�U�(���F�<_<ޚ�S�a\�px/B�s�W�I�[	���������W���)��Qb����'�GB�J4,��l��<��6�V1��ZŖ�v]��,���v����>����s�(�~UG��&N��_!��<�N]�m�]M�M9*���D�3�$s��5��<���������d8�:9��k���0A�̣Ua�\0�*JۊN�@�"�oGWy-�}P
�=�o��_%i3� D��B�v{�EA@>�e���ҫ��z�(j�
�0�O���/3A�RDh�Yy���>�WH2Xs��ڃ�g�����/�c'(N
e��8�W����3��ux�װ�&���@�l�~�Y��Zu�Z�\��=X>���1���c���k�h��)*z_�&	wp哌���O`�mvE���=�����m�U,̏���hޅc����]𦶻��\*����0�k��wmaNҾ�CN|k��:8+�V���^�.�w���m�
�~��J[�vV���7I!���	�X P�����.��e�oe6�]�)'�"�o�!a���c@]�%��B��v|F��<�������W�^�섞@\��z5�H&���D�CDzzϵ����r%��ڸ�������Z}�UU���kn~�����9����'G;]M��ܑݥ�e����Y2LF��Nd��������J��ے�F��+ו�G���R�X1�@��\. ��5־�����M��}��mY�ۉJ��`��4Z&ͷ9�!9�OuF���c���h��!>DT�K���I�����m�J!{�	�vA�*�bϖ�uX���<�y��!Ӷ��ӌ̰mc.X��;���z#VF�
y��9�N���k��}A)z���F�ZH2�
�L�<�>�U�`"��Z�a[��.1�����!%Os%K@�K�L�my\~-�P9
���6�:q��1��d��3%�d��<������z&>M�������������gaH�r���9���n��@ۼ^�_�#�$if9�]�A|¤�t)KX��*�m=���w9Lba����d�I����϶C���AH7*i8(j`Mz�E9/8������:��[�ī2d+F��0�y�(I001T�x��Y�7`��ds�&��Ø�[���	,Ag�:��K6�u4_��� c���f{���&�b@*����y�$��]g��z�0[���F��a	!E��� �V�B�`\_�:����g�p�GgA	p�w@m���E.3]�j��������9º�bG�=��U)J�(�t{��
@�P:��ꔒ���%B�3�=3 rXȫȇ[H��|[G�6���f�D��QEϰU�Iﳿ�R�{hAd�����kL��:�� ����6�$Ia?.�@���"��4�9ۣ���u�9����=��[��g&J̌@Z��q^(��*QI�Z#>�����i\V���ӂ�Q���=�e������gv�����K_1��3b�����-c�{s�]�L��,>��&0~�T߬H�CU�Z6�M��G{*Bd�ԃYz��j��[����r�7�R,�g�SlX��sG�1٨���6j�:}���3���wƽw��7U�c$�:�EI2ų&E��x�ea�⏴�	�z�|�"�<�&;�ī/�ꦍo/�EM�cSn\����0�Q�d�~��܇+��=U��3&���M7Ƒcо-��S00��E�9����~���r�m�Y+$Bd���:��UB����F�p�p,7���H4.}j�|9+��,q�q��e��^���1��-@�	��/qm+��W��b�oc[ui!R�3��{�A_�zz�B�I����)�Vw���Ï!o0�Ī���KC�2��bŎ�F�LS%�VmɸRRP/�$n�rZ����cӛ���<�W�I���CI|d�g�,�|2���?L�p�-[5�JZ���k�}�t��|��d=z&���c�sX1k��u���}��п�i����1G~w�Ï���6��\u��}V[H�99D��&�S�O�>�Bp=�4�d�|x[l����W� �i�L���g��5��P+�7�)��!N{@�h��7ݎ��Y\Ǻ�[�
�)LQ��rו����s�����q>4�I2�A����V���jA���F���[9�39#�k\��,��˯����y,4��Kl�?�D�&|�>@!�3z�n�Q��I��8�+�
E<�ӿ!6K���xϒt��씽(ױ��_��>���� B�I0�Pv�Yj)�>�<����"�4e���u�R��~N�W|�)��ԫ��j7+3����b}�	 ��p�9�t5nu'�b���`�Ai�DbB�Td/�h�ʄ���2'�q��|8M:9�Q��#aO��BavT�*��_���L���ٻ�̽����6p��u��s���e!�$N��@>���&[����'��t�y�^X���S�Ӟ[T��m��~�s�qk2��^��i��J��� �].Yc�}iz:�HK�#eCFA�䒳�֝�����j�i�]��	&ݏ#^���&}cHoQ!�j�e:
���J���w�0�B�U_p�Q���WOyND�'|/�V%I~#�A]�u�f�6�h$"�B"�����G��i<F����p1t
�E�/[�=x�l"�Jua�Z���bF�oȽIb� �'�Ο��<'pj`�Cq�\�	9�ƑT�J2�8�ZV�!�)�1�si
�̓3���Bf�&�G���$u��^��q����Tg�yi�*`|����)!����
&A�6�v�����vA��T����i+�V�G)z�ߐ�e����aO�=K�U��`����Ȏ���֠�m�}pm���5!�g�:i�p����.����L?~�@��^s���%D#���v�Gb�F|�ʙ�|N�r�|ppY7C�c���
��1U�8�z\/�\�C-���pvm��L˕��֬�Gؿr|nhF	��p�G���k�<�� d%��x7`j�ssV	��Q������9jO��(�1����q��o�/�#p��k���O�P����%�W�9Aތ�� :�2G�ۇ��T� �vҢMN���wD[��~-��M��T�}�>����Q�_(O��}�!at�*�Yj�J�0�V;���V��l��mt؇��
�o��V���Uȩ!�06 )��Q0���
�0��E�U	���y�D���Q���?=��8D�$Z��m�#�Ө9M��Ee�:u:�ݻr�.G�S�X�k'\~0^�^�����x��9�BK R�������E:bĶ5g8�r�6t)	2D~�X�M�漱�ڳ�TJ���-up�-o�E�}���'|L�U�P/�8Rn�<뱂O�[ɳXh����;4���`��"��	`_4�#����%I��W(�����F����?�Q�dBhA.(��8p�o^ɜ���$:۬I�WX�N�K=��^�@k���1]��D,*Q�(���֋�M.ؑ(�#M�#s�'��
[8X��Y������/(	Fh��P+3O��_��_�V:%/n��;}�%���nÜ�e�A:_y6DH�@��=��Ғ�_1���NI���Y� Y������見��\�C�@S��E�O� (�&hʱ5�l�K���w3z�ם0&��v��
|��N�ӌ�j���j�]2e9�b fd%��y��aX�F�A�K��ʰ?�����!I��d$�Q!��ݫ�g���X�e���x'w�ƍ���ĉ�s���Ǐ���8�z�F�O�u�s���ފ�p�)����9��J��#����)᪵��Kk���q����t��2�#���{�r�I�h�2�+�JE�  ��9�B�8�cX��*��2'�ʉp���n��UIv^�����L�8>r�v��D)_�]Tl~��|j2@/�z����o�D��l��v~!m$�ߒ�qgy��z6��b��{s�c�s����?���Y�.yH�0:'tg�M�gf�}P�L`�D"�� �so�g�ZTZ�x~��d�*�b5��HNKqݬ���\�Dj$����V}���-ͧzoC�#8�E�����b���B�΁>�!�嬯�����Aq1_0T�
R1�m�T�K�,aA�p�θRQC]��-RD�[��d��WT��x�����ɠ�u��p�ž����7T��3��)�
ֆSRROM����,7s_up���0R&-�;��i̿�������'U� �)mC�{��#�����t
yj�Y��#7�eA�:�H�TB�O=t]����Y �6�ؼpi����
5��mwV��lɹ	�q�\��G�t��|Q��p�=+1��}ܢ|��+/�ۃrr.���L�s�������{��ğ��J/��x�b�F6�!����F�!B��蝳
����h�������x&�V�I=%]���0�J��-�<�%#��2�'0��&-9mA�&S�7��<p"?6�!u�wm��`�h�LVe{}i�� 4dk��'D� !��Fmu�0�5'㥌)����F7�tSOUI"��=�����;ZJ]`��Èe6AN��Dvg^oW��
��d����;�D�g�d=�o��v7rxu'J"��9�WS�f��_ȋ�6��`O�ՀM[�ˏ_�I���tR7���"��8}�6���?��=��9MP���V�k{n��q�Y?�B��(k�?eb`"ζd�^|;qX�ʧ>O��<5u� �k�|(�*&����LZ�ݺs��
���_6۷wVY�q����F��ëX�>G��z�}0�}�ά�9ݮ1f�
��GR��bBlyI��D�X�Y�������ˮert�94?Xw�#������@�5c�ɡ���,���sb�S-�ROj��c|]���Y{��в�Z���l�=��;*��2���#�B��
(B��C��d�_�9��>O��(����C���9L*�f��:n�<�����y;��}-�&���HY����"
����{�3���h����N�ik�/�\��������)���]��z�p��6��a�=�5��6����z�к��M���p�_��\�4�>\q��P_���~�3�7�WH=��eh��q��y������kط��=������	<qu���/��������7H���"E���L%�����ޮ�	/n�f.�� R8<Z))&:Q�9-/��L���di*�a{��N�L_ì��*��"��x^����Ҧ%ٻ��1���~y8H���h�ns��iD�o�E��j�f��������dt4w�bb��j۠�s�x��	�˫+��m�:�JB���d�E&��Af7-4v�XwOh��z�i��q�ES-
�mh�G������Rz*�V{��e��S��T�>
�hT��'(�p\;���&%�8��.�%�N�ߧG?�|]L2Gq,�t2�j��*��o�98G���/<ML(�����o�֛��H��$m�h��=4"4Z���=�d~9MM�	i3��%����o��2u�HFF�*QH>�T���2��Z�/��f��p��d+�db�u߸	D8����"v2�+AFI]�H��7�1����P.��Bt�Q)fo����p���6_���0����NO�+��j����Cv��~)��

tnɌ�K2P�F���sѺ0��h�J�<�mቿ����սA�t7. ���70��税����G�@u}@s���'��1�;AI��R��Ϲq��Z e�x52���w��R�5�f��_��ު�j/���Ϛ��-��>���g��T�x�~��ȳ�"�tb}����F�� � BI�F�1`s�%��P�?:���]�;��6*���t]��R�춘`�9��:[X_�q3��;��Y�t|UoT?���6g|z߈�aˤ'���ǚd���Vy���cQ�*�Fǜ��P��cq�s�^Y2V��s�yY���N�:�ӿ}�0UqCv]���C>W���}�t�i��#����8�<#�U�_�����l�����~�b`6��Qҷ��n$����ZnM���֧G�����j����7��Y�[	f���VB���@>���W2����$"�{���u�R����e�8h%��wT�� Z�qA[m�����/��` '����	>��d(�l/,h�4�
JQ ���.��_��TI5�b5L�(4���0���qKcF�N �a+{��O��o>pa8�V�n��f�`-����J�(N{V�u,�D�`f���[��r9T�{q��ğ2�N�m`\�3�G�zZǳ��a�N���!�t{3������>��PuT[;�ܴ�����oVT���1�̇���Zwp�!G��D]0֎����%��x$ȠG5y�_����A��3K(���K}�i�Z���R;2{��Z+��öUZ�����~|�&���@�mVD7>��:tb�bEQ��\t���LGWz���q�������˒m�$ t��'e]�	�:"�`9E����W2��%2�Ӈ�|�v�;
���ǘ;*a�AaS��:.�A�26��"f��CS2����܉��kkV�}��:�9�Q��6YOO����F�YA	���D�/�Gk�3%�a��)U��iG%^'n�F`��"Z��A���J�AکX\��V1PUYS��/
�B�BU�x�����A�%z��ͨ��H&����+%?N�R�
Z�S��^�`dE����7[b�4pX�z���ĨP�(��]�S��$����$���A��B���'�iKP�~[w�К5
T�D���0��z:\��Zc8�
V��$m��{�!X��ښ�/�rB��l���pv� &���B����U6K�(�2ƸNB��D�� =,����&'h�R�$���c���*����F��қ$�G+o�J��=d�?	
�j\ᾘ�u=��6ݩk�/���n����`��iz�I�B৻I�-)�m�u˃�Qg�?E�p{�z�w�a�HIQƷ�š۴���ݡ�[��\�E/�XmI5u+؅������)5,l��bX[��C�v-;�*��� es���l��+v����d	��`L9���ٯX��+��t���M+�� Pp���3��)܆��-��=���!|�=D��+|u�U� ����?MP�X�~S�#�<$w��	n�nF,⍇Uo(��(r� �͉�]쑭!��z뺺Wki�� ���\�]PΥy��V���揬���pXo�!�m���NI#*/t����(RO	�.߃�F?e�к�q���L�.����i* ��5��p�X�#9VW�?�Ŗ2c.4gx9?Pg����:��\��:N��]z�m<,�+��"B׀��:� ��F�	�㙹<2+8�}1�'�B=��c�x�ې�Mk�����"'۸�	�����k�/�'��Ƣ��_A\2�Ϧ9�όm��L����LZ��|6`8��]ؕ�&�׿��F�Ɔl5E�<'�>�ނ��"�#��`X���Iwc����ī�vf����ZM
`$#���f��9��e¯���/�c��]%�N�G�n�0��D�.-��>����i]���߅d��n�p�F@�!8�Ӏԛu_�'Y�5o<<,5��LV��$�v�;��q��hK,^��2cѕ���Q�!\_N �v3�"pH$I��]oWS�ϴ��w�h$łvv*|�Cna	-�xZ�s	��E}yW��c��C��;'���g����$ڏ�Co~� ����O+y@����lo<�,�'g'��y��e�A�!C��x���{D�)ɍ�.k�i[�,����n[�34�-S%a*�6�^�V�%��+:�i�G��<����!�C����F�մ�}8�01/=g=�ST�n6�]ʻ�w�f��j��K��!�:P�_5���c���B��m���t�
�Q<��$C������h��e�3a�,�Çm/��~���̾6b�f��DG3��G�#�m����/h8� '��t��7â�3�I�Cc��?��������X��u�"D�`8}�B��X��J��������>�Ra�p��r6A���D,�_)��@����C,����A��iӘ3Uo:���e>N��g<ҟ��֨?C*���t�|w��
z��\ޒ3�u�#�k6���Y-�?6f�V{�v��� 2����$U�d(?��Љ^�b�1�2_):h� \���`�D�U����Ţ�-���t-�Uo&��3�K�b�͔��h�~N�J=�`���ĕ�|��r�jU�����qM�׿Ձ\܃=��E���f����R#�y��Ѿ]-���T�vĨl����D�Hf��}�6Y�覯x�jLk�h��o�5�I��j��l�E�/��:b�Yl@����%l�-y<�R��,	1+e��h��ZFe��j�;�Ai%��'!������@1'^�r�Y��·	oB-�W�:N�
�(���b�5c��#��OU��j�����FTR7��a�}��-�N����F�{��Um2�F��?�G�]�B�;�{��f➒�zdȎ[nK��!�G�O\'���!�@^�\N��t�r#���띃���xJ�W�+�2�b-�=�x� I����-��y��헏s)�w~�������u�j+�{!J͉<%���ҡ�A�'�(*��\7��	k홧� ���m�Q����#{R����7�cJz�����×�~SWewGta������8g	������4��'�lޘ���j*)G�B�`��Qз����?=��9��������n-���j�|��ܮ�5+B�T���;���$���P�ߣh猡E���\��`�*Tw샒ros�)�#.�\Čk�h���E���~W�爮�H��@���d�?�����3���qkXO���V�$��{�kL�M���r;��(UK?8��lM�;n��k�4��"��	�!#��������[�r��0������U�U��ҏ*#��ާ��b�ળ/���B������ZȐ�@Yt�JDݖ���j�H��>�k�]�,aX�3��g������ͪ�,gu5�ag�����w�򜳞_0ޮ�W�FT3*��{�kq�14-$��v"�#�T
6�h�5����Q�Zj�XD<@%=r�n��z���,�İ��{ԧ̆o>[�,i,a�ئ*z�T�4:�����v��9r�5B���Pʮ~��N��D׳�զQx8���\2�E����"���́�~t<n��m׹8������hAN�*1��4/�k�AM [b22_Cz*s.0��(�Z_0z2�/z���B���Y�P�bLve���&�ȧ@�c�j^6!
-�A�!%��i�a��/���i�_w�өFW��{���*4���e8�
�*�"�]�.��S�Z���^W��[2����ɋ`������jP�B����G7�U8
ւ�'�<�I�!�v/%Ԟ��ٲMq��٘pO��Q����S��;�de�����xG|b"��m_}5�cF����u5@-������{�Ѫ�]5U�/�W�%˶��Ǩ�y*���f-�QR��ͯa2�,jd�}=�j�^��\G��ބ9��3D�U^��!�!�?�q���Y����aO��`D�O'���JD��/~�ZQo|?��W}fQ٤׮,�0��B)�IM�u�����:An���?Y��`'��~�-`�cm��G��΍�9�{����t�Sm�%�$Ni�h�rH<����@E4�~���6�O��f��w�F1�*8�wU��M�М|�:8ϥ���d�
v��!��&���6�e�!���c+4���ѤU�EW$�h���(�h�&�Ma��&?��x��B��U���?9��t��/c'�������é-��������	K��?��L�����xde��2`0$�T�HׯtП���r�I�t������RD����~_��[f�����dS#�E��Bh��*�P���j�Mn��'�`��E��A륇􈝎�$���J����Ĵ�n���u1z_e��2^�3�;J������W�x����Զ{|O���T�Zh�A�n�3�Or��C��Az��~�����iF���*w�!۪�7��� ����P=[���D�ڦi�/�һ��������T�~��
Ќ1o�(u*���i�DŌ�l@G
)EL����� E�c�-1��O퓾��j=��dNe�l�*���у�`[F4���j|aߵEz���kG,_�=¼�.�;[s5�e`��6�yR��2j�*TXr/�h����;59�/2gIZ�-����{�t�c0��W�g:������/��9�����8��K҈5��"��I%�@��z��K[�d�+�=Z����n�4Ke0�T��E�����]���w�G>���jC��s�ج`;�~z6�Ӡ֠W\�ɺG*�&��b�����Z(�j��\�E�ۙ�U�!$}��v���4��U�@�H�S>�F����[�4_�#�@�IY�=����@i���M��<4��TyO�b�)P�W+k�~�3���c�3����9�2&�d���\+g�fp�"�Q�����L��"����2���0m�ki��<G6Z�jϊ��nDx i~B�d�w��i,�o7^��N7]��k�J���0����W���x�#�\�t�0m8=C�
}ec��<�`���%�V�(�;�7�j,��kCa���<n|H�w�x�^�r;<�;����>Z{���3��&�ؓ��+̛f��ߡ���@��U�
�+d��i����1�R�W��W�U�
hYY�dXe�Y[�/yc������g۪�u�=P�,ޮ���L���sO�Uq�7lyW��FO�y	K�i��8�=QW&0�c!~oS]�Q�0���vR�U��^~��z�F}'J�'<k�u�}^��J�~9��`���D�)^�*�-�^�<��r�,�	Ў�%�o���������Y!�	�LWrup_jG�c�n2��f��V2��������//h��@S#~�mp���C}H�4:����n��J��%M"�g�����
?���f�υ����.ǭ#R�nO��2���P]��^��h���ª��g�}��Df�)�c�4X�����4��ܧ��3�T��q��]����/h�r//Y+�@,l�췯�Xa��C0���v�m{Z]�4���v� �y��t����]V��=�f$(�@S��D3�H͔�~p.@�xW���8&��L�S�k?�T7ɢ�g7��4Ձ�S>�Cb�r�%0����Q�y�I=N:�C��+�z1C�OLAR�p�L���h�>�%X�W�F�ep9#�ݹ�#�u�|����T��g�)��3�ssVx����z��L���Tff�p�t�q�zu<��~�S�Tb�w�{}g����S�Mb]�rY���p��������]L������KpFw
�!�`�N�EIG��E���i��-�[rJ��P7#+�{�RoI����?.''>�R&�w��7�^p�[��
���� �����;��NW84�'ڹ�,4n�B��+��p&��2��5���R�8����c^��z�kG>���@P����ۡ�,����^��zP�o8�G�#�?󆗉w��٘���O�[��)
Ld�`��@sD�<4�8#n㞑Qn���
hR���p?�Wq��e��h���O����z9�0쬈B�ä=��,4^�G*�wIY{�4%|���M��8)�4)�h8c,}%����aҟ���M�X�*-򂇇T-�����:<�3�=;[v}�X���*�MƠ��yg�$��nj-Y&<�T���_!�
rS���%<����P��ߵ
����Î���A0�/����Sࣅ�}16]���NU����I-��^�Ruu��:;���.H|��^�ţ�d�J��Cڸ�cf�c�>�l��m{e�g�KUP��]����q�d,$�PꞂ�<U~�nXXz�5�ID$��b�}j�s�ge~��ɵ�E�L����:�
K5��2A������G��sIf���۵��a��G6�Z��'�I&E*�ׯ�sF<��k�~u��z��]�l@������%!�jE����Q�)�T֪�������=�̈́�a��	^83���=�ZC�����[�����s�ԗ�����<$,۠[�����pu�#��z��5��T��ڭjn�CKm���|,���C&�s�i��M7f����?)X��Y��i��(�*�{*V���'98N�+Vh�[bFX�a$]]� �L�KBTl��b�gj*bJ08�EepeN��J�v+�On�/¾$��⾫�o��Ԇ�u C�$�C�̝{S�>YC���� %����E��\����LjW�.[	b�;_�qJ	�_^����"X��o(|�{p���&��8.����޴� ���^-����1t�j�J���.t�O�x����	�f�i�Ԡ9��U7��4f4���嬢^pE�?$4?�=Oݲ�+5b�;��4OND#���y[C�+9�?���J*k�mҹ?��D�=�smdLe��&�h�c�w���i�Oo w��p���tKXpԞ�X��/m��a9����C+7�ܗ�\n\�I�x��.���4��N�R��m�ݩ�n��Z����@�1�l�_���!φ�5��~p�MT�;��d�D!���ڙ�^,�Al"c���	�	�J_Ϸn�~\jA�Q.���v���!����� X��ݷUĠ���+�{�s��J����Y���b����1۝�vL;�*١[��wJ��R��JmM|�<0�2�������7!�����WtT\豎��QR��XZ���ۯ��5~p�q��.�ڢ٩e�G�p?;'��̜ͧ�lT�ϋ�v�=���9��a��i"B��f���� EoF����_f,%!'��%�,Vʍ��<(�o�y����U�����D9��V��Ϋ�y;�j��� ���} �����o��iGVUZu3��� �p��e�����\{I�#�m �<tV�套�����Xbp�~��J))�hw7�2���0I��^V������q��'���6�=9_s��*8DZ	>4> ����pS�g+2쳀��lԓ�zH���>Q�PО�+'?�b%	/�����y�;:���g�3U����v���J�(�|L�4LL���ɽ��\=<�����@��,Y���I���!�]��h<��8<��ɓ+�/?�	3N2P�S���EՍL�%�p*�ļJ;��G�a��}����� 66�6n��J���f>�!Z�`T�A������BcT�*��u�ww�o��-P�*�d�ųD���""�g�����$�Yl7V���!�W����˓�&#�D��f�ָ�^:�6t����_���{욇Q6�ZtU�o:�g��VC�|�gr�[��J`҆�N�rD�N+�*يǓ'���i���G�\���?́�{�*+�ԏ`�V�g��
p�x��s��� �_�I�d����I�T�8�FgHРo��8"���^��,Պ���r�Gz�2H!N��U8AkS�Щ��Aۢ�(�m�"o��xNJ��`8��P�EP-�����C@Y:�a�N���'��c��Gx!�|�?�>AJO��+�\��6jְ��.S�C򡵖E�����JB�_h7��D#�����!C^��6�I���CC)�t!4��F@�D#��a�hri��c�[�b�<�x��P{1]��7J�C������
��%P$�1-��K$����:��	^�>��P�"�k��C���Q:Xz�!��f�є�I�J>�f��͍�l1Z���;�ߤ�� �a�5な5�PnB�`X�EI�<�1 ��v�ȅx����'=�D����\^�G�z��h[�Hn%R���^&x�Ƭ	r�
�k�#�jpW�9��Ęe!�m`�=é;�S��<��L��H�jh}ľ\�%�^�hQ��Gj�J�q_��jg䮲�:�w�v-�EN��.���VҖ�*ߍk����\\����$�Q�sW[}X�6���[q�*N̫��N�-�ε�����<0�%��Á�	��@t95�0cέ���}�=ϐ3&<C�V�j�)9�;�p�� �_5D�O#���!Ӱ�JwWF�cÞE|p�X�ukl�x?�ߌҀ<��]"2<�!�6[���8K��3�S��P🡥����/:�e{;1���^Z�sk_7��|H_�y�~ۡ�����$ٍvp:mYwr��q"4�+��>p��h���1'����{��ԟ��%��"���� �҈\gkMѳ�� a����=4T��ߩ����q��wU���c��Ư�]��`�9h�[���<_ޔҞF޹�%s�J(�#Nq����� [X�DD/+�k�c2s��)��e��d9�j>kؾ����;��� ��X<��i
Q&[2p99c�:�x�<��@_��3�!�K�C�Cݦ]�J���4�������]�|�E�dP�Nm~�Q��{�\�*s�0�`�6mW\��)ߔ�°ͭ"�@$�r����U�&I	=���i�e]U��a�o�����, �BM�KMG��FH�XB=}"�4�8�9,�Ga}j�%����0,3���T�4N%`��5{�0� n0���s�B��B��qV��7]$�I��dG��!��u6n&tL��I�o�x@i��ٜ��i:��~�pҳ�r��/i#&���א�Sq&�j�z͌F&�'��0���	;�E�u��0��>i+i�$����15� �j:�'�i�W
n�Ts�q[ˤc�c�(*�qd�`��9�E-<quf���k����je��t5����'��B�TDv�� S5� ;@R@�/�*����
R͕����
�}��U[��kmkέ�U��q
��z�i�k_xƉ;�~_�T�묤�=��R��Y_���o�m'���ʍ�텈 ������x)��:�KJ�z�AD��U&�Vp�(�´�0�J�La7J$$�pRg��7:}�1�،�G�Գ�ZOL��%�"j+5�Oq��-�D�#�!�B�V�=@�G�Y�1R0�A@�ɳ�����	�%[�y�X~�퉻ؒTa1\�<1]$R��\�'����:�՗�<�&� 3_�*� ���  ��O��VJ������iP�`	ϗ�>
�����X�	��k��Р�+���-�FV��?��|m�֤�^�Afo�8t\M$��������
E���IXn�L2z�[�uR��̷a�(u,��V����L��}������S�<�Ie�/��Z�9�y(�|��	�REުX���`X��B�zI��l�\(C� �&������46�]�B�����{�o�����Cd�h�w��Y�4�aن��P����2c����g������єrL�+��t؆ *E+��1Gs���~�v��aȲ�O;V�ا��E��A$��a�I����Z`���.�����
a���Qj�A��2���GQ�Gװ��8�܄%'���7 nWia[Q7�����$+��:��'x���oo��(q�����TT�KM�P���S�
@�_��i�k�{��'��	�^�(��S�ɪy�|�L�DK�N�u�{"=|9�jk����j�s���'ټKNϠE~��D
v��]�p��U}_�&u�=�VNX�\�r�`>7�B�x6ؒ���(Ȗ�Y�ެ�Q��nw��ǈ��t��ۿ'�7�sF�aVN�q+ͤ]�ƕ����X3���-~(l��x�,-��7�D�E�	m�Á�!e�(���B���Z�v<ia,+�	 &��ۨ������v/ e���*�ֹ�Ą��8Z N!S[��}q?n�P�����JL#[�����6��w�M�)���2Yz'R���L��b���f�����'��SBͩ���p�LQu^@����\+��RMZsw�&�n��G����K�{q�%��� ����r��$�`DQ�]���$
����p
�i��Ek�=^Y❣�i�i�G�	��/��݂�o��ef4y)>�U	�6_0(��M]o��[5U c�@�I��'���7�M8P�����R����ia�sGS�CԢ��ن���4a̎�'>H�S��p�qc��0�!9V:m�p�A����P�h�Uגq�^���,Q��¿,T ��>�5*�QL��]uyw�x]�S���8���#�*�xn����zNY�����m׭݋J�]�B�q_د�"y�'�_;���@�2�x'&��+��$ᇏ�>�&巼�x�ʉ�h<p��mw��=�f�N��^�Q��h��f�G�P�急�]��f�}���i)x)�G�<�̯����k�#�fl�R��v�l����wJ����]�[F�0h��E�G�v�#�/9lg��I���p�h��7�rѼFP���Ҍ���4y����ȷZk����Q����������撲�ڊ6�Xzu�� QMM��Y�b�CL���_7��.�cn��6ljP-]2���MgP����7��K�e�
�[l	��8�|O��ckvE��YՒ�;�ք�_�c�$�=��ś"`�o�����bd��c�'ඃʶ嶹��8z��H�H�X��fM�t˴�gEvg���!���䛴�P�?H'��LܘZ��:@���u|�i�U�k�G`KLx�N����!/3d>8��C�h�O�K]�'K�|&�Gvv�8=�'�g�qTQ��d/���'�S&�'2�.>�B����%��S�i�?�n��ɭ���۝�@�?��^j@3�  �m���K7!��r3̦���`Rra'%���Yuӥ�s7��O�D�<�A܇����	.!sX5�����֙�7=�����F��B����Z�`����\0lm��Q��>Q����w 8&5��OB�c|�񟅪Pn%k����Z��UM���ɢ�|ƾ-k"���^z���7���X�!/�#��K;���A!�����ٵ��3��9d��T��7p]p����)v�δY�$j���a�a�b!�"p�լ�QF���%�v�n�]�G,6g����2>{��:��fp��\�Լ��Ohx�q}ɗ��Yvh�3��h$��w~�yYe�ȒU(�uQ�'�&ҧ��=������9%������5����b�i�J��͏]��&;��D�5~w���8�v5�P��fH&(��]�ږ���ӈ�-���k4 ?2j�Ns��a���M��X.A�/�`w4�z��R�p3�� �bԷ�ƺ�Ei��{��&���VY�T�������-Sk��?盆�ev��Y�
�֡���xџR:�C�}u��X�jˬ]ਾ�z%wB&?�_�m
�zS.���E�Iq�&��� �$���(-����kZ��4��ݜ|��|\�m�5�a�� ��;����'�Oz����Y=.��J�Wܓ��qPW�c��\>�qƃ$8$��àQ�jM2�l�-5 ������W�g@R[��R�r�;n��Mg��.�T��]~4�m�V�6N h�W4zH��@��܅p%��,�yR�����īE������M%=�.��%k��j-�i��>l �a�<�{����[�Os�����i����q��Dx1��RD)�T�.ϴz�?��7�3iO��H�@��\�Hk�)�d�dV���Y;0@����$��I���%����S,'?,Ñ�Rf?̀�i��6�3 8��<d&'K%��"��p;�B�]�����(�B�����D�<w�&[d}�s'��a��9 �8_�E&\��6%:)BҀ�L�'�dz��I�X�S��"��Ky��HY~.�rN�fHb�9��L�6u��������쓯F���$t� v�G|��,�����uH��<u8U�� d�_��� t�H�m{���x�އ���PI�%*�#�b�Ft���d.�#v`AI��
��oz�Sq�^Fo�Z��U���.�xK�s��5�$�4�MNy0�ռ�.�������j���[p`�������W�S��/+�z!n����xB
���b��;�(+���O7(��R)U�<�;t47�f����[=PK��LR���3�M��e��ƚ�Lp���Tݠ8~.
'�Y����%L�0��\5���
�e�Nn��:�c�����~���aw��7����= �[���HmrR񶰥�O�Q�+|����wX�i���|cr/���Bṣ���h���&'�C���b�8�?4��.	�V��绅�j���'�o���u��Ot�%<cf�4k�uN��简�'ia�}�7pX�	� B�������jM������C~B�����ס3��[�jw�� U<ݙi�5��
�m����UV[��nY����5�T�-�e�{RҨZ:���3����2�žnR�ӹ�"1���>���g1B��Ƹb*=dܖ�Cq��k����+����@���.Ef_�.,w���(�g�:*�!�C��J��i��R�Q��I�	�j�l6�����c�������qQ5K���gk����_N@�L��U�AiM����͔|�?��j���d���Nݢ���D\��� ���m����t۩sQ�)k��K�����W�'��x���s�fd2a�`~29�h�1��t���Ⱦ�`&���R	Xk�ָ�%��1F����؇XF�e!�-�ן��f�J6	�A�5�![�'�;�zHR�"�����f���jSe���K�r«�����e�\hTC�m�B1.��kU��<�8P��Ë��C7����/�B��WR��ܸ:ݙ梟�7T�[8i���e+U�A\j1��W�5�졒O=��*���{5��2��%F��@6m_����q8��QE�����ģA�O�m�<ʪ˛�h��WďqĠx�B�ޮ��g�d���<,���l驟GbC��v����4���/q��'r�2�7�,���!�k�󩔮�ږ�.��&�� �f2,R���ۏ�Y���b�yZg-M��2�`�_���(��x!�����+5�~ZT�$�7ܩ�əl�r�J5��K_��ܜ,ԃ�@���G�m�Mzf4?��}".ۗ�ҏ�'7gj�`S��>>	�$�hv�,1"�s��|��q�+K���#�1�e���1r�w&���'"��R`�7�L�ţ��#�H�{�� xf�0Ϗ�����F�q��=�Yp���j��i="�T֫�-�{Aˇ}M�[9���]ங�y�\-m�U�"s|�JK�Z���	���=z��t�L�Wat,�Sʬ�^����(�N,�@�M�-��g����t�C���[�X�K�n\Z���D~N�K��V 0����� D8��5�L�V�ʝ2;Ε^�ݢ�8�b��S.�f匞#ytE���Q���=�̦���D����Ű{�ܥX@��0�����P�ӆw��Ad�J,ǲzQ ���?��a���ѓ-�F%�PDf�V��e'f4�t���`g��oZ(\�}�ߥd�Gɢ�	UTZTa��3x�
.&p!<���^s�=������
;�B����i?���n�+�`[B�Q�3rh�㧧3�d����e�"RV~�,���\B5�V�� p� ��4�p7n�1%A#�̉���v��}��'�U��y��k��$T�h�����5�q;��m�p�v0�1�&���u3Š:���Cٗ� �	wD������p-��ȑ$	Ԩ9ʇ~�1�]�� S����ɕ�> z��V��+��T+��1�=S��{�~`��]�#	l�0bCa��{������8~4&���ܘ^\/�6Z�Vv*O�s�O�s#���'��>���/~��\�]�'e�8���8T�L b%S���6����mUFh\2���[�H�szw=*ٱ����(W�u'ZPLL<��o3=8�#�w}x��A	�ˀ���K���GW�/��)�A��a�jCAOލ�Ty�m�v|��[����%���#�89E����E1X�25߷lP��z�����h�m��Na��~�gU�N�ॡ������Zj����ɑ��m���R/N{�$�`�frh]��� k쑁~�7������"��IUq'�ʻ��
/��I���B=H"euտg�������4W�@}c)�jt�Vt ���QT�m!�(jǏ�o%*�PU
��`�P~�
��N`<x�'�{e}8L6ۦ�̖]��+	K��6�;+@no������)�-E��z�3lل�a�e���@9=����"hK��g�� ���Lґ�T���5Fq�eLO)��qĐ��rm�p�� Wr�8)4�^����q$���f��J 1����c�o
s��m�nΡ�sx1�,������~�`�$-���ڡP�&^�1]���Բ��>�6j�,�� �$i)
��lKp�,��S34���f$���;��l�����{�Ռ!h��j>w��ٸ���M`�s�'�g�Iw� `�s��b^�h-�G�]�}N_��5<�8,� ��G����#4lo4���1}a�;D7)d��h�[W�ܡ.��"kal������<M��ژ�+9yY4��y���E-�>:pN�^��c(��i{yZy]=�(E�<9�G�$U�����?��yV�_'�B�"|�f@���l��V*�VڍW�(�&�>}ƌ*��_�y�y��Ӑ4NPףΦc�������ߔ)�Hڅ��^����_�7��G�Jb�ԈP�4v���E*\�Ş��ꂘ���6$�%~X�����f5�Q�.�T� �l�hǀJcY6�b��a��#���G!�<����[��b"�����L� ��o���:����<�c��	]���x
���v*tl7ˊ.�tV��4@�¦�.D��zc2Y$��)��Ĉ��@�*��Uf@l��VZ��h�b<#��N�ۛ	"�����Ǭ8�j���"tpjc5?p0b<��a�l�DҒX�E}U�������s;��&z55t�\ew�U����Go<���SS&'��D�&�D!���j슩j�ƑD�ە>���;y��U���I<ɉxásb�+�(��}d�;-�94J9�@¨�*�@V������c>���S�K���5��ݜ�a�v��0S,:����5@�|U4�%U�o=8!'��h�ߧ5}��/�([�؜	���Ć���/�[C���8���'	T�|�����F\M�Ci��
gC� � & { T�[K���'��?�idu���E�A?�#�ȏ���Mϭp����Y��f�<�6ؽC8D��z]P0�j��P�K�炘���K0U������<�T�n�F��'F��@d��Q�������_1Ł��vhGY4��C|"im��:�$]�}����w�WԮ1RSe�%r"�<VU�^m�W�B�l;��v�Ӛ+%���b�����C^P��MpM$l�P(����i��-�0�b3u�h_�;�ޖ�8�s��x�l�/��X��)G��:CF�P���Tt�0+=��j��6�J�}<(���8!r�GW�ßN"�L���,Zv�ۛ����\P�Ǐm������T
�Y.|���56���P+E��IJm�GM�-
R]�_3���X"��GK�|���j�ɦ�n|A��3���7fYqC�+�(�b�7uS����=�*#h����}����'Q��@S��ݰ+�G�	�qMd~ �zr�=q�܋��0^JR����Z�*�u�������ɴ�8�޼�I�]�!�	ӳ���)�n�G��B5P�m����zU�
F�*��v���	r�$����L��
��i�j	�J�__C�<�A���p��O68��B������kUc=�>��D��=�$i�h�A.\p��N�8�}�O�(0%#�Y�lֶR����T�N�xY����W�p�{2��O�AM6Ju{M�W;g%�O��&b��5`;,w'�f���E�PI2�i�]z����\���$
+ӳXJ��2���܎��(*HZ��8��6j����/�Ƚ:&��$��?H��5�����qƙ�+la�b�=�<���U�������7�ؙ2�8�31ɞ&�`��B��u'���R�"�V�DRB̅ 2��ͅ8Δ')�=5X�M��4��d�9d���E���h}v��Uu떔'�֦����/�v<]P�V&�y�K���5��yT�/��#������c)B���
C��R�.�����	��-��~����~n���//�DyTf��Q�őiαҊ׉�U?`�Y�?tiն|��r��ǿ���im
c����0�ҒWc��1�Xj����e�Cb/�̢a�ً�'���xw�y��%�����s�i�H'B��^,�͆�_厖i��b>�cg� j0H�tal�tO�$:@��O_8�,��mgH ��!�N����@�)��' ����O:N)�^K�t�h#Tr�z1Qm	
��U?��ւ;*g�P`�/���V�Z�����,�P<<v��Ѯ󾜒miy�2;֖��j��p��ݚ�����},Ǝ��������@������N��^!����C�|���+aD�ل�[i;�.g����۹�4	\v�8�"��_s1l�\�ѿc�{����p�@���\r�j�-�x����~����iӝ�;��B�ɷ[�j�*ӳ�޲L��p���Ǭ���It0���[��y�7��|w��J���cqna`t%��,u��MG�.Y5fy
v�:wK�k���W�]�cn��T$���mҭ��[��6D�Y���'�/��q*:��O�x�䒞�-0p?G�/��y��6��t��+����\V���ZuA�Ͷ)��
Ȓ}�v��Jv젘���B�����HPo_<����W���K+�P�kdU,H%��)r}	��ߵi$@���>�{���`�5�(l��#VyS<3%m-�`��G�LG6�����}'��T�¶ܖ������4��Wyk\�V:�W�=�X���`�&�<�D0-�)t����-{��T$O�B��֦xI��y�u�\�W}�S�㹳�y�� Hp�祙�J{��(��tu_Ifd�B�ƽi7�����goOK'Cq��0�~���r�jط�1_��;k��σxp�_+�-���-0����h2cv�i$+�t�C���h#��Q7��N��2�L��%�����s��q�߉�ݹߓ>�yY]aJFX(:�`��؆{�4"�;G�@�4��|¦���Z]�>��a��.�!��=��N9�:���7�q0t$?��	�u�z��}/~�n��/�:���~Ł
�n���S9�I^�.қ0��S��aKr�7��Pi>���M���MT��|�KW�k��jʓ��R)K����Z�ڋ�ݩܶ�^c��vCӗ�W���/�U�:������&g�1��4�|�*C"w�y;�N��ז[]H��a��/�b�m��#f��&*V��pV�
�[̞t)��ZG��|��s�o ���^F�)1�@�r.�ň��� ���d+f��D)�^��8Z��ʎx���������z'�G��5=:u�м�C�rqG���Y����^��N=�	\����K2Pͩ�j��bc�v�9��/s'q�J�`��Mz�i1���j���M93m����CHt}�O�������&��mf>U�g��V�n4��2v��ﱎ\poF�0����b��)�)�W(dc�;h���.�j��g���DT�9ފ����B٠�ZU����5Vȅ
���}/e;r8l_&1����i��df0�/���D�.;Q����y����-l �UɄD)��Z��v-#	�4۞��g�7��!Fꈚ��D ���rbZ�Ӑt&���|�|-F���U�Rs��d�gӮ6,�r����Cǘ۵6���&
�������a�{�j+0�;����E�W|��+���"L�iu'�.���O
������qv��1�x7E��c��<�u0A٢�|GHXn!m{�l�Jb�ski�#��@hC�{*�ɪ��S�ہ�0�����J���97{�4TH��bva(6=�U95�8.�˴�&]~�#h��������� �MV�
����
��D~!�P��[�ړ<�Z���9b�g�lh�dɘ�:i���`MM]�T�2��TL5N	��S���ύ-H�����KJ�޲0J���&��|��p�.�4�Ό����#�q��l��K_ANϘ�3��:�`a5w���/�{�ˡg�3����M�Eՠ(��݄5x�a�9�&�:mS��̤HO��I+q����iU��KP~NV���bN�]�����
fX�B+�IVqL
!}�������H��ⵚ}w����h��v ��B8�B��]j�s%�@�r)S~'_��7����Ҁ'�Y�B�'�,Щ����א*�*3�M�w�M홓�ϚEn�f-XX7@�U.��ٴH���Y6~���C,��8���4SR����J`x��T����Ѹ���goWW!�&j�$X�ǟe�v]<4�N�1�0�4�M��^�[ J�B�\k&��0��,j��� ���+�����D��2�xc�7��6�F�6��Q�T���fTN9�r����:_�0=��zf�g\E؊�ݔ����[��-lr~c�ƲO�8)�?6������},9w��/�Ǘz�<�0x���A1 ��+P�kF��W�<V�%�6� �Y�c�_��i��� *��K ��h;.��v�ߝC�f\e��Qj3����h˯ok^�p����q��;��S�ϞDA$C58�y��E����x��P�?��O�&�ܸ�P��!,>���%�����/�Ͳ�?��I�ۇ�Ұ>Ój���S?2fl�T4����>H˖r:�zV3�s!�Uy�����# $m���)�\�/�x>����*~�-tГx�2������u)9wC�b��8\�/���8�uh6�[J�I�F-|5\�)C�J����H)r.��B/꾆Y��'@8~I\�H�f[�.o����]��ah��Q*&`8���ф�	_��1�,��y^d$g��63���hN��ʧ^�c	�5��s�GnH��r�+���`��F=�tf��/�u����37�O����/N�%W�2Ah��I��F�M�����NR虅Y7y���TCh�my����c��NS2�V�@C�I4+2�vg_���p��+i����fyP8�ˡ�R%�*6~X��[��-���C� 1v���D�-�-|�%"��Q��p�e�;�&�!!-L�}��OV��q�fs;�դ�Ghaqa��6�)�؆���&��7���d����
y_m�p�~��zCG��Ǔi��	r"��<~�Ø��hfdQg�%h��zv�����/�C�/�������D �؇��Wء���� ���/^���4��Ъ-�)����J%�����K2���~CYl���{��+����0��~D���a0~�֘���$���z�D<&�b!gL�A�	1Y�vr����^C�!�:K�7��EF�ɉE�A$C���$�q�8�'S,	��|$�%�/R�4`����%�"�T�Ab��{�KԱ����݂����=��_;�#��?�+Q[1 �N*�J�Q��G��4o�3)� Km`o�S^K}D�-����Q�6Q�� �� T��ү&F�bZ������Y�j�ʢ�����<�1�Ϧjb; ���Eo!K�\�w.�MB0j� �Z��O�6k�*^x��� "��}-��&;�t�Wk1b���Gr�=���_�`�w�k*rs^̭��ti��oQ���Z�C䃲����Q�"f�$la�#�Yy�:�V�efn׃"��1<"��_Z#�Z��1��K9���5J�ҙq}y��� 4�:��U1R������q�M~$߮�W�-"*�k�}N*�o�l!��I��D���Q6��`0=F�#$N�(?��Dw'�v�lY��
;<�<����|�';�Ktњ�8l����:cf}��`�n�T�6!pR�NOj�d/�H�1tI)�e-N�wʦ�����T��$[Q�:침R���?��*f�N�54*v#����=�v{��K�:���^Ƥ�T�)�!�&N�݆R]�*������r K�3���z���`^5@/��*'
W�1�1�R�*�>�H�;â�O�����y��?��5#s���h�L�Q�͚�d٦�M�r�\�I�7ʀ�R���vDn����q���|����Jc�Q����i7:xy�q��Dx=�p��%G�AiˑZ�"j�)]�5C�����K���}�����Gmd����{fL(�_'��̉�á���ܦ��ۈb�Yh����݀�'i!�i sd��.ll���wl-�&3K63�a�!>�Dd^u�`�TuG3Z�����e�
G����:�u�������k~s� ��3�E�V�O�T��R�Ѵ�!d��w�"��X
��`bW�)��j���l��ú�#埤l^ �*h����A|�m������eϬ�`� h�g#����/�����=���p���J`�9�B�=�r����E�X��Cl���*�����-��Ѓϩ4�
���e��!X�M-#.l)�6,��l�˔Vi�Џ�)d��B/�T�!Q���V5KwU*�o��!f�}��߃T�rv=7�͈c�Q�_�s�-�6%��xˢ�j0��#[�=�\�Uc�%}�N��(�����c����?&���q���ܛ{x
��k�Htĸa!&(���eZ� �l*�1���o��d��T�E�V�@涻a~;х����^�wS_0K0�x����d�� �p#X:��(y������{��(���c�������
 �1iP/��$"��qV��a� ����PK��G��d�I=������"�@+Y��Q��;�@ǣ�RC?���}��Qle�{����w-w�(�w�ӻ�_`%�>�M�f��G葃�"ɪl+�@j�y��De���،�X#V��C!�uĨ��ϋqL)�_��x᥁D+���	ӿ��ft_��4e��:e�Ew�K6')���<�y.���CI��D�dDղش+M�����ӵ-�~��! H�J���y�?�P/4IE�4���#�dC����a]��N���E"=<����,Cz� �Yi*ijp���;Fl�!�8�G�Y{&p,F7��1��6w���3�P�$�uʕ~��,�8�x�D}��h���nڠg&���B������">�@�Eb�4֔s� ����3%.ȷK�tA2"5Ңa4�bxH��%���JGv����@���|������q��y�X��LɢC���Of���7��e�0�2"bTH���~��>	9dR S[y�A������FE["�cΕ?؄Ȕ�'��o�z�2ozNkf�-ä�=I�l�w�e��s��L�O��\��y,�5���l�CI�VPz[A~3l.��b�1�ޱW����n
���Dt��&�jl՛��
��U�M����˱Ó',XM`�J� ���+E���3d`�x+�`Y�3�D����RH�ٞ�бD���C�#y��lD��.>4x@`���϶��	Kl�6{�{��Sv�_ͫj������wnfBz�����������:�q�座�c���(�}�_1`� LW�r"��`'��o[-,c�����s��,~�P+����}�����������%\�a68ژ�\q�;j�x��]�l��Ļ/L��y[�	�#��)��R2�/��1rJVv�ڙQkX�]%��� �|t��r��㰎縵 �8�����!ݼ-��� &'߹�8���˄�KT���&되���=�-�9�0~_$�Z�r,��F����P��%[蚴ԇ�j����a����0p9^OQ�1y���s�n7�i�y���xZlӡ|�\K�q����8�f��#CQ��Y�j�/�{x��eag�j�uU���fB#�bāM�>�0�	�+r
��4���)n���F|9̇��#:�MAA�~��2��G�~������tUgr��8-�W���g��%�+��ڳ�#Gۗ��2QTxb?��������>���1�h�m;~��^9b��������[�R�4<�V �,��< !��M��)Z���M�L�pW����~�Iƾ9Z#r��oak̈?;jHE�f��֊�ﳧ~׮'��O�k�6�b#�é\��H!��3i��� .݄�<���ƳJlu�Lɖ{�Y0�����XC����)؞��c%F<I�17�����y0U�S���q�+�f4����R��`�(}d�P�J�YmeQ���a���0Z�D�{d3-�'N��`ؐ�Is˶f���]H�5f�剩+�������u��l),/��~��޳|�|�5K����v;�R9+Sn8GgX�#��I��d�#*;(�����Is��Wq!A���.b����ffi���,�U�ŷs$��W���r+J�\PD��zs�y�ӕV���UP���(�Z���MIb�n���*[���o#6��A=^\d�6+���ȎU'�O�rЉź�/�(����d��S���N�Jf\����ڴ4B&>��r^��$�4���Ot>�;&�>��Z֎6[���v�Tn�u�.V�F����a|QߘA,u��Y��c+~�g��������4#wq� ���)#�hƳ�����lO\�_���\eN�Zg�yɥ�zğ��|�G�vNmQ
5%Al�y�2l�({'͕96�������
��W�U������O+f.�K,s4)��hl�&ǒ���uݢD�Z���.L��O�0�Si�P�ם�v��zTF���W*�2o�Ρ^�L,A��,��^�W��.spqN9������N����πD=�jJ������i^GP���R� C��ܦ<�&�k��ٺ�������\��0����ph3��0p~}��p�xyz5�)�z�Y�����\�XM�[�#m(o�gK�"�rZ��{D�������ez�m$9�X�n�{�/���<DC.��C*ҳ]�< WŰ)4��_��d�p�o�k�+�z�ϲ��~��ط�(NfEI��E+Bk������d�b{��U���S�?����<q�������s���1�.����XC�^�1.����B�h�
^0k)�Ƿ�(����3���4�FX�^ ��#țx��]�7|�q�2��L*Au���K�<����9����S~���d��Q�&�5y���0��vg�<�܅�"��M\| �1�%ꡉ��u �ʄ.��ܿ������5�D��L����{�3�R�qt��Sj�[��b&n׾��@$�8�M� -�a��L׸ �Gz�a�e���sO|$s�Ϙ�I�yߝUV��V���|�y�S��>��m�s$��8�&Z�O~O�j�� �c+ˀ���_PV�P�q��\�ܘ�_{�3MX��OUcJef�J4�Af�a؛[+'���M�8��_&b8����K%�jZ�G2�'�a�/���k��*,~����%�����K��c/j��*�G��.MM�T[E�;3�45"�`�v�F�d���1�DCf���g�5_��B�+B׻�coքL`J���m�8K�c_��U��J�I��%��5K/��׉Y������MևhBYʪ��/���B��9�/Y�r���
w漪���ԠѤmS$�"z�� R9(c�:�����M��r���c���y)X�\�u����߻eal�:|�>����a���}��hۚ�Y-�'}0��5��t��2B�f�A�����a36�[R�c���Qk¨6��߮pbN��"y�,u=�e�ڴ���b����e���*���ldw�h���f���@>]��,���M>����͝��KS�`o5���#�w+��N��E��
kkp4}?o�Z�ZP*vlmۘW�UfV�����7`�5)i:j�,�{�]���}�3y��*�g����Gұ3�c�?��]�Ep<1N����L/} �=etm�p�(��	;�/�4�y$�S;�s=��P���y|3��0�i�$b;IŠ�z ��翊ޓ�+��H���P�x �?�������4���� s{k62��^�&�q\�)f�nk��UnzY�%l�R\���&�vR(4 �F��Q�{hP�!"P��Hov"�~!�Yi�+�PH�V�����%Y�G���$��~�yP�v7�pB�6!b�R ���?��<�������D~��,�K`
ڂT�����lY�.x�v`���(2zLz��
"��b���o��*��K����{�<��gG�g�.�)����v�XZ� �Y��Ng/R��.y>�%�#��;3?$�2�������(>�����LyH�R����Ŧ��N/�����փbi� ���4���Z���=����B⟝����l�G�j�4Qm^�&0؃NB��f�Z�8����Ep��N�!B��.�'����Q ��0S��N��:��Q/��wgKw�_�����ģ��ʥ}n8�i.���Gsdc�2��=!1�/\���Y���U��%��0�zV(v��L���nt1Ɵ?νpj�yM[�AA�����.�+��`�R��N<9���9o%�9K�a,�̾�(�B�~wW�̦ky�H'1����n�?5���t��=����-�@)׬d[�%�����P�n�bY)��������n���FX��v�����:0��8�bz��'�����p��c?�k���U�Z���C�J�__�1�/�3�����ޖҝ���+�I�*HB�h(a�NĿ����V56�؜TV�D6^��4k)GG��=���'&�U�?PA�m���s!�H����5]Нf���ģj�߇	*߁�G�8yD�)�W�X �{�����#��޶�f,]�'�[��e3����$�G\�Ƅ��wW��HU?�g,(�vXD����Rx=��b:��M�J��d�ژ�k_� /�B"�����!��!���y�+���F3���.Ư�GQW*�6��>��:�(�� 1�)�)�V���O��"g�?���J���y7�S�lH9�6�Kz�� %-y��͂��^���K�T����W&?U��b��+j�����}�M��ׂ`Do���D��ա;xZ�Fqͅ���6��!V/[�����\eTEg}�kċ�r�~��S��ԉ�`݄@�e�u޾�K�G������b�W9`��r/~"-���Gfao�������Qw�Q��e��^ѧ1��O�܄�7P��kw�UB/�etm�[���jk��Z���%���L��?`��þr쉄��N^�H��w���M9�J(Ē~�;��=Y��&� J V|��>\�`m�ԑ��y����x>��t�ʋ��s/I�U�-n��I6�)��oY�O�7�F~��51�5��h�C�٪F�
�+4��S��әp�`[�u��R��*$}4o	���H�mP,�]��v��U����sh�-�??u2�� OY�h�� �3��
V��v$2��Q�nր.@�0z������>?��(iSG��&��a���}`�������d��$��1m1��i��WK���^vcƮ�zV��W/<P'��:l��@�eKl���LH��R�9�Q0�e���e3�fЉB��ƏS�`��f�44:�`ܨ=�p�@jzCa���%hm8]Ų�g�7�jy05fj,��O��)�G��,�m��,�ӠnkD����p9�6���Zbԙ�� hR �W�kN4����DԎ�*�F�����(xz@6px�%��qƣ�ؚ�!<zGhf여A2l� �Om�����Ҏwa	ŉP�2v�2�f~���4xle4�BKm ����%VH5��R�c��>���nЫ��� �A����Cմ��`X�v�\7[%�h�y��o�$v��l;������#	������[�.��{�R��C��7�,5�w��&Q�Ҩb���KK[XN�By��2��Q���vB��db���ȩ��}�<(��r��ĮVE����Hh�τQIJ��h*�ǅ{�ޅP�F�eXt"]��1��1+�<��Q��Ǚ�c��\�S�4�bV>%C���i[6�3��fO�'�9�y��#��A�X�o2��מ.�VӚO7�;�ng���hB7L;[m�0k�{�W��"8��2�*l7��IW�#�<�B��Wђ�	vO��_�qTm�r��!Vm�I���X�mj�~e����M�5�)R����A9SO�d��O7?ɽ��S@ �U�Y�D ȗ��m�M�ĥ��+D#dW7����Q�h�	�����D�io���c������
��5.bk�f��ի�i�-�`�v: mi�/~����|a�j�\����tY����#G��3�P�R�o�
vO�7�O�j�Q�Nx|Xɏ�n�_�IR�o�/���#��`�HPg?2��ˑ(��j࡛K�R������ Z�K�V��d�	ۡ��H-�O�6��:î���l���E��'+��g��������pFgJ>�O���c.��C=������K:ʂ����+y�^�y�Ë�����%_�v�O���8H3�1�FK����-K*哯�����(��bH�<B�����-�0G�@��&:&�l���_���(IǼ���g�
�n��ω��p����۹1M�˝�gr���`�=w<βBe��;�X2@�Gay����jȪڡ�4��/��������G,dD�;ӀN~��n� �ii�UAQJ������e���S�`�U�H�<��2~��X�"G��c�I�� E�;�5�����L�o�D`�w�u$��ZU���������Ok�#\=�2	O�6���-�N����C��a�j74��\�-&*�ڳ�<��Q�6��%,:�85��0�6�V�akv�*h��Q�m���#�!�7C�0�%EC��l�hwwsgò�@���rVQ��^=��_�פ��jl�̔��A��f"M7�`T�o�2�E����^.(�X�ۮ�m�d`�{�`�
�����sg�~=�ob�kz�ja���zk�?��U�)����]!�DB�<����i!ϝ�w��v����z��L�[��a�mS8������w��b3�l��P~�ﭖeU��HJ�)~�L �s��)�������������54�mq٦����(8�9��,2��k]4@������nI{�y���+=H1��W�[ b�'^�s���;��A��K�F����b^�t3�p�������?mKD�~q�d�q�юu�|Ɯ<J\ʹ�Q�G�����jqUe����JU(��>c3h�	g��B�\A~�[v�̃2'�ED�/�=Ï�eRp�?J�%l�����.)���	0����?��[��^�-u_|'7��
U��J�Ԩ���p��+�_��%�d��ג{$煴�έj����q���&Rf�i9"�Ԟ�f��}��
V���}��4��E��MFJ��`eK���e��7���3���ѥL�c�`�g��p(�D�`V����Ժ�V�[5�n�Fb�~e%eW���G������c���Y ��P���)E�Ag��C�� ב�O��s�9bj7�(V��.X��S�9|!��q���u��`�d.�V$��2?�NE�����"�����	���1
��䙢Kk���/W7��ܗ5_�l�|2��Wg���-aX�����O��m�q�ux�J$�']+��|�Dj��@�J����3ċ������б�D�g=�?��Lc�(���z#"O�dƾoN��Iy��7ca���9���f�|1� },;Bv�w�S�qP�I�"�A}�&;����Y#+�7�΃�	%Mkõ�����cf����.��n;P��M=�v�l��4����}{���!���j�Oy���%)�=gM�K�ߵ�X8�7�G�[�W;��I���I.;m�#��f����YzWeKf%��O/���.1�֕.��y$S��^��PI
d��^�r�:�D�<ҝ-�0�a��w�LiA����,��튧��+��2�9{r��%�ɞp��C�7U���Zj|,��+��4��314�b��4�Z��=�@�Z�ؐ#z��2�����κ��q�N��[ꆠզ>f�f	�C�~�e	��̓1�4m���j#R-��=���-ӷTm�X�0��q�11�^�;�C��W�b�+�Q������pOt�nk@j�Z?�I�^WPzR��u�%µA��J��;oR��>}׍��_�SS�<L"�-��*�OrL��̣�4�JM/|� �#��w&"�p^�B�i��{�-�HO$���~�4��K&0t�
���{dRZ� )�v���N��+��١=Y��!�ِ�?4�TGd�ĝp^8u�{�n����͡v��ar<���srC��M?�4YkJl�돠͂�]j�Ȯ��E�G�o�u#4Xi�n-$�N>�̞�\Qz��l#UϽ�a��������u?��`\���L<Q��{}�Fux:E%�>Q� �^)��7��S���hy/��N�tag�%�X�ؘ���9�#��mDgib:69�O�l��b�9n���T��|=�qf�b{K�eG��ƴ�H�@9�폸�_7��y�T�(�(���&��_9JҊT�Q�a�p�ʩq�[�����-���;�	I��9 	��}�p�W�X��l�$ ���`�>:6\��ʣSн�/$�2��_��q>PZaxk��5`�0�k���K�|@O��mw���:�w�)�S0ްk�W<�������`��a[d�i���pW��m.
���\bZ��hq��/�'�߄m�[i���:@���7CCX��e5q�c.!f#�n���[�"�\��UH����$��)"�K�� *����;�Et���T)�����BHb᠀�X����n',��ɞ,㥛.�/5.>k����΢�H�Ol
�%cu�grK���8~S0��8IZ���L���埰��&�)P�#4E�6�O�����m��#�w�zh���j�wU�<]�ż�8�>Cl㗩u��,�"I��׶e$W��N-�҅S������q?��>n�$b���Po�`5o��U��s��`�R��i���7D���ޑ�����seΓ4�/*��{�x�0ʋO[ͥQC���B�z��_�\��DF�fef�[�*2�i�JK����9^����	�\��f-����](.?	6}1^�h,� ���k	O��h�!]ΰ�ă=W+; #��q�묞H�2���O��c}��Zٌ��}'�F��i�'��]M{�� )�y�C�o� d&�W���gh_?PD��V�#�,/M� ��iAg�FN�F�8a*+�y��$�2���d��q��vb	,�)�#����}y'YP>�h�6�����F*G�n@H6�^7�ɴ��Φ'ݚ=�����흂U�W�\A�� �1̌� >vܼ`RT{�+P��{!�^��f�z%�r.-�<֥��3����p���o�YKT�rexzv+ꝑ��7!S�/nm���^��5�h�ý��\*���D�mC��1�'5�ӄ9i�xD�	����|�'Mż�V��+��{X*��B���J"����*��3X���6^([l/8��<�ť@�<U�S٠�,�p��k��r2Σ��p7?�K\a��4�n]��tb��PE(|]���)K:�Zx��"��3Y��7���/��%㣺�B�4���]m���O�2\if���gž�8cf�� ynac�b�(�H�x7���\K�s��n��b�G�_׋�bd�K��Zԣ�ǩM��
�f���_	~���,[5�m~"3D�䳪XnsS�^�73BP!�B��`j7Y@)+������uh�<~��i���-bsR\"�<曍8N�������(�;��80ϕu,���2�.<,�ɸ���.�=�r�2�m���$iI���z�G�z��5�L���f}�L6���+���7VZ�}X�����R�y��y�TT�֓���Ԡ�q�\h��~��E�����[���[�<����c�D�m�qq3����D�����w{Z��>����'㐇Q����bD&z���KJ�8��H�[�؜��@��C5B�:8f�Ӫjh#F<7vf���M�6}�Ks-�=S)�An0���sDm��D
���_��I����C�_�g����	S���d���?xB�7��n7Kw �����̖04��G��0_ꩋ�j�E������_r�������=���L} �B�X�[���ؔ�AZVWw*̡yG�������?�5@.`�������®ڿ��i-���ue�GQ%.���7�Z���7�d�3����Z%Η��q�5�>�|{wz[_�s;�&�5�8r��=��t�?tI�O@]�Y����`�>e�F��-�F���(��Ѣ^�Z��#�?�צ�XR��cK;tg�Kr�}	�����n�z92� �A���Ĭ)�x��G���J3hx9ʣ`(j�c�୒�>^��r� �;��B�f����[{����x�5������WTA �x�.�Q�RE�0iw�ӄ���4�U�k��eDٯh�j�λ=J���Vl���x޺�MP�_�[̐G�Z�|�2�-�n��k��X��L�j�B��IF�Ƃ+�$���h�*kg1��:wZ�62m�'�!t$񅢠	My�Ճ�r��B�r�o���`���dlX��V?�c��O��Ƴvz�	�B��ؼ���B��f�Ο�Il�Bǡ����߻#�X��|���^��ո��.�#0ʏPi��t�Q��p�ݶt�/�v@�{�K�����\�S 1xG�9q^8���R)��I�4��lΚ��ZEY���p'3Ý%0��	q�cW�'�Kg���b�EY��Z#�MؤaD�}H'V���wK��$�M����=�Q�\��L�s�<}E�P˥T�j���^p�w���W�%�9k�/�����V�~�?�z+eZh�E����v!4�2��Qk��K�D��'+�!�[	 �Fi7�-�5��^\���&9[�)0��-�kq:����g�I���H�dF!�J��t�Xޑy�y�P�>C<�:��/��\����H��k-�?\씫��WL$��f���x�L��C�qH�=�)v/lT�W�3B�e���~���_�6���� (��;$���C�A
z
G���5+��F�c������AG�hlL{#�?楶����gL�^��@SVr)�*rK��y+&��Α���Gp�\h����r*��(��V	�;�GԜ˜ �.�V`n�et)u#&�]�{�W�;�L\��=ƳS��w:p���P�x/�*�ہކ"��ݛc���f^�_�j؞�CR0Їl�7�\ �+=��)��]bK��'��#W�iVa柁չ�l�2��l�@f�gĮ͂��ԭA�B�1�h�Ɏ�a��#�se�(0A�/`�bV>���^{�Кo�����O�[��a�e����N�tW�g�b��ϧ%3n�!z
��ڥ���I��Q��6�.Kv]��fw?�b�̮��Ġ��\����Sn7)�Rk�zғmu�u��:j��W�ܚ@��bO�혗�_
��%-Ԕ<�>�,�m��$@�9������Z�b�{9�-�
Q��L�𛖈$�̊���?�Y���+��q{��@�4������s�dtٌH����+`�)w-�Z��B0��6��.�E���[�);Jx�rDޛ�Z^�bڇ[r7��tݲ<Zj+�*vPэpo�ǎ�U���)�)���Y��>YQM�Jۿ8�-c�)uD��W����I��,�j�`�9���"�w,@�lKL�Lqj��nH����?*l��d8�|W�<�ۃ͂��ե�Hr��v<�8S����[�>J���l<��}�l��7tS���%<�)��5��+�.�o-����K�J��[��E#sI΃L��5����u����&S+�)�4��L"w���zVe�s�
����H�;�����?�hD'ڂLRe��HϾQ�7�6/9%O��i^���"Tz�)�t�}�����m�'��XMP�����W(��&+7%S����	w�2:�a��/X�X�h�i��]���X��0n��}�ǣD��*��,f���`�������>_�T�Z&@�:M�V䴀���8K���Q�j�(sr3ܞ\�r?\�t�/ٻg 1���9[�s6h�9�-�U�{��(q@�0����Ή�JT2KμR��c��^���v`OH�5��NN��Nj�%;��)Д���,OoC+p���d����w�Y�YY��	 �J��ƙ�,�]�W�A�p�T �.y�懏Jhi����:�SC��<
���f�I�6���bh��>m&���]���ôY?獃
}���L��,����N�U̖�E4ꉒ��z�A#�3U�$|�k�X�����25��k�Mx.��e�a��8q�.��_�a�Q� �J��r�����q��M��u*p_��Dg�jj�%C��;*F��.j�`�j�J�ն-uVz�Jp����B7R�������t�蔇#%B��=��.Z��^g���z�9bw1(N��������m��q��2��kds���c,���"l��,�<���/�P��V>�i���c)k>�l
���lxg�Q��YE��WH�����ε:��w�T�7z3(l���7�nqfDeU�L�a�ע1$zrR�'e��Y�n�g�;Ucs᏾���B[�G'��w� ���]�X"��/M��{�����:� +��_�B�m�e(���5aɲ�w��:��G�H������Vu��05f	�P����9��77����'�IŴS]"1,��L�`��Y���co6��<�
�,�)l�10�V�a�<����Y �T�5bc��@��4�����n�>�3��j��m�Z�-a ÷I����	ZIFH	�V*���dg���ԯx��¢cQ�'��8����74Ǹ����FE���,D�f�Ķ+���T鋺C�8����(�D5�$�Zk��{���� )F�m3��}m7�Sh0�~�y>ˊ
�J�ԘZ/�P9?�z�
`,4I�(a�,ʸ{s��*	���Ue�?�r/����#�b���r~��т�l�(���A�Q]�������Ӌ��o���X�R&Id�>r��;��XL¤�5��|�@}z�'ί�=���6&��)ګ�6͢�6kS����mE����_� (��8��#f$;�z�T�A��0^YR�U*h�Z>fU���g��Ր!)�(C`��L��Y��$��&Ep�&U��µժ�$�6����I�ku��yn0�k%eq`Tݩ��TX���nF濞��Z�m�|�Q� V�"����2?�k-j)�Wޜx�_��9�d8��̱��7R"n,�hy^�J�X���jZ_��v�V��,��N���-�Iuo�^~l뇇��K���Dh�t�_�(�	��J+�\ʇ�c��9�4Rqό��i���j�γ�1���$G􈸛u[�/�}kǡY�q�}M�D?;j�(�M�i;��������y�J���=N$�WZ�����QYIIC 2�h
V�o�?сEg+߈�n�G����G�Xɬ���PF�q�9��҄iO��y� �W:%P�����Ʈ����aID�7�pG&�H�b�.�3�rA�#���$/�"�����"�#Oo]����KK����HܩF8���i�V)3��������DS6دj��;^��M�X�0��ͦ�c'�ХL8Of�a|�da�����W�+[X�EO�%Z׶�l����V�K�nxYQ���M���Y�ju�N�0��r1�[6�ëf0�_��}�wK�T�n���B�\�����JKD���ޡ�K�����*�o�6%���޽�\Ch��І��gM)f�s�-Sa�%�ժZ���"�+1�0V"����D��V�:��to&�'P0�����.��+(!���	#�{^��Yc�b���׉��(����22���O�����L,�Weġt��v65�`P>��6�8�o9c����Np�)cSl|bX�0-�����7��q74辕#�'vg���M5��l��c�I�L����|��)7��]�X��[	Y�B�s��]���;�"����r$���*EBR�o�sy�L���
��r��>�ϕj���>�R�� �������"LH����T�I��r��dI"��J�n-!���6��h�%�����.�f�+������JH��1���0�.�,wn�CYD����.�zk�F`�M`R�i(�&��jtA�^�Nr�����0�V�Ďg�"�`P����ˢwY��o�I���0Y7�拉��v�@�ng����J�\�,�F��Dʶ=�w���H�_g4�E� .q�^,`����?�H�z���n�o�
0��;D���c��FX<�R��Ǚf�*�ܤl/9G�C�۝U�8#��I������(�h��vsXS����Ir�p���3XP�V��:��0U�=f��D+$�ǃ*�{�e��*��K+�7I�(6)G��il^˱�1�G�%/�!��O$��t�O��f8�f>KV�LS^�|�4�,��׼.s7҄c��j��𕯏��_���2f�� n_�N��0���}�-X򫚵h�ڧ���U�-Iy�J�hE�/��lc�(�s�`��� �Zt.���Q�3B�S�l�q(�g�Т��� A��`��������ځ$8A��8���d:��c\�"���c�?zg��n���s�����8J���U�Ty���ʸ�f�(��R�ӵ�٭�����28�.���=�
Î�{��2G��q�f<߇}�e�%I����KD�g����Eo�CF��Q恕w�s2��r9�V��@�=��R����(^�����]�O�ӓ��b�o��oE��r�4g�XW�/�W��؎��여"W�$�`�*f�_)�\[G~�B�Y�>���%���o�ȡ䋒vXp��hg����j�؇2�ZUm�~Hm�<�\Z�DGyzSOlU�M����ᶀ?�$���0n����J��>4�tlA��q]~�3�Sn�w��:DT�0�`Yc�$�Tգ��O364 �T(��e��|~[.]DO'�W�ظ�oǘ�r6t�Ӫ?��?�i#⁳A����)����r�TSU�� ��Ɜ��)�`�$�GLp�Ȉ�?�v��2g�kj����"���ƙUg�9���|9=!OA(�b)x�������0̋jZY��%K$ܸe�g�m��v�g�	�D�+�00>���ƥU�,��k��9pi����f�2?�/`�o\`{�k�8�Z_H	�\�<�5�(��椙㿐��>r�6Gn�<Z���Ӧ )T��2�O�\hcRUy�$�!��G\����si�ɢ��}��4'I0`/*TǬn�Z�!�Uj�����Jg�APv':"�o��d�n270Sy���J���no	E��׀�57����rA��2ޅY�Fm*\��@D�SF��Z����s�x�d�N�M��R,�����@���l`�#7G��wr1$*�H�����H��c��&k��=b+���G����:b��i§�σ�x]p�C�b(a?����{��pZ _LI	�[��H(�T7m���ƪ���p�<\��
���a�H��t��]����� ��A��0�:iW{[�$|��9.�÷���m���B� {�� 8�CrF��_�c=r��U;;����*�B,ڍ���60���)��.%�yyA�
�$A���8�ˋ�Y�b���$�(_|	u��s����y�w��&�u�
����H؈�J���&����sQ9���:|yOeJ��f*���?�~�lIR�V�I��W�v�V���8c��xJ�S�>�Ҥ�d@���I����k�B�_���;"r��rz9���<��ٚj�d2�i�U�96�{��}�ǌ�����g8Y�G R����K��Rtl6�_�������E�Y
�=����d78�rdW�ԉp�h�=\b�����w�C]����Iy��,�g�`�N�����K�� �N��������>+G������dУѳ[�H����2�a�,�	7n����ע���̛�]���l��I�(��ԏ6�`�ո7Ћ�d�1M¼R��T�U�H����5G�� T��j��W h5�����E�@��t�L����b��52�!�&��(�}�w(�R�����X_�bT�e�_���Ƨ�ZF]�h$�O�������	=���	������iX��N������}����Sŉ����e6���z5�زkߍ�ۄq�!��	5U=պ�-�AcA%�7ϙ����+�wh�dm� ]�������M�� �Q�^���tea����Q,ό.c��]I���J����a�����k�"�#5W�~�hIu�Ms*�Us�٤Q5�a��OB�'��6��� ����%Q1H��~NUfߡC&�"GK��ThN��;��T��A��Z�*�r5��'吝��uq��J�xS͏h�"����grQЈzGqۻfU5WV`	���U]�1$�b�ݫ������g����R?�Y˲ڱM�Z:܀�ɭR,h��yԟ}�"��zm�E�Q����K��2m������*���ƚ�}�,x����x�f�i�Ci�Ϡ`	2+�.�_�hԘΖ��'��y�����9��$��>�^����]|}�#>�J���8I
���W��'	�	)��t1D���A�ݻk	����<�4ِ�[��Nl�B�`���MA�V��τ�p��3p8�e;Z�>N�U!gL��򣄏�B��m��xR]��JHR���;����6��f��/ �64�@�j�$d���]�m-���6�ڮ�}�����x]jRd�\�T���[ߣ���GԮ�I�1k]L�i�T�j��G}������hd_�"��}�=�6���L��%U���߁�m���7f�����-�t�l��� `I$����96F��>Ah�,��}U����Km�ψ@l�	���-lD�7���4 �֔�UI/`��oc77u]���gr8B�^��f���~��y��ߞU�0ň�'l���U~����1{��>{���LX]�&�@���-j���6w�3��t�^<�<������>oD�F�%b>Ŧq�e�AT	�M
s~�@<V�E��Ґtu
��!�J���u���t7����t�.| ѣ��I��|���޶*0�{Qp��ɖL��@#b��3�aRLULFF)y<2�w�w
Q+�
��.���ɵ{Q��&TA5|�Y�{�d�R�����d!|zJ�4����u�z�
����y��~j���{2�0t�ZOg�!X�E�u����zP������4��Z�ЙK!Ϟ��J�2��J�'I|�F<��/�])c��