��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��mX�Պ�$��0�s�zw�
h���4���.}�mA��,�d��e�%:�}�+��H������u����]�jז��S[�"Qc���qiS�kDj`�����7�5G��Ξ@�,��]��!��_9�������{�d�[��o`�}������M@Rć�4�S%H�^��m �Qc�Pg��B�A��L��Ek�����W�٫�]�#�@5�=�1��灵�١}�N���>�s���#�yF�� �A���h�H�: �^x1�Ts$t%���*%�:��*Ry�r=F��ѿ�ʭnh�Q�����ݬ	kѯ=�,�ԥU!�C�i8"�)���ŷ{��at��IK;�fJkM���ǘ���:ͩ�
�pb!�v�X��O|�9�T�5��GGl��G�F{2����cWp�)J�	�~x��y;eM��jh�4�Ĝ6l^��]
�;7,�7�Wi�>=j�{��V�m�" �t��4�O��9�R@8����[I�mj?� �)��Z��N'��ſ^o_=�l����n�9�n*���-7M}GvC�D~��9AOlj�bg���>���T��U�)��	���Yl���Ro߭X+��%Z�Q���Z�_�n�T�	lh���9��j�/��b�|�B�=�m?F &��#�%/1v%2!_���y�/��~�X�A	�3�g/(kTܱ RE,]4<0Nг:v�7���m�Ӧ<|O�ϺX2c�q)̎;����,�+�|מ������_t������Ujx�/)<�"���F����}�E��h�|7����ג�jah%<���C����J:<V�D�Pry�m�H��ў�'��7L�V`�#��J쇈 �X�Y����ѭ�� �)�!����:c|���9�}3a1�^�r�8"Vz��&��!+�b%mE��sfe4�K�Q�ZJ���T�'V��h/B<Y�A��|������Ҭ���m�gHa#���9	=������j�e{�x`�
)�o��+�A-RfŅzP���$�Lٻ�0少J��1^̽���S����:�˵�Si�f��bF�(�M�#���b̢�΀:7�����ek%�
�$���1��B����ş>k"p\���,��Z�'����m�yG�ÛIjݭ'7M�� g�K��&��;��f���n�kC�B
ϯkHై��>9�Qr�'����)�~v����Pʓp����`I�O���=*����(X��ٜ4�0TX��,��C���+&8����EA�� �"L����<c��Ԝ�7>8�G��7f<��?�U](<�g�n���U1!�3[�0cUq��]�w���J،5��r5��V��~�PRO�Vi����~��w�b�I�Ҫ�a��/��F�?<�9Ԁ���q�ʉI"�x�5�KZ�"��a��a���I��(	�s�)�+�|"�.z�O��mu��~u�n��A�@�2��q+P-�22�ʇ?u��f�
�XW��&���G
0˨ơL����62�F�_���A{���E�`������ܱ�9���_Ʌ�B��<ƀ�
Jn�.t�n���Z�>e���B���i���]'�gbB�e��al� b��:_�o�boBwMs�?A	H�������y�lW�Z���@������"�<a�����Ǵ���k���)�=��zL\׬����S��ky�V�o�N#KV%�&E��d���N���ZF�iD��/YދrQ6)e��fRҤd��U�Wk�MU��2	B%�+�Jq�(h?4{g����|L0���_�rt?�~(�=q�&� QJ���~N7�8�8��ZńW�ވk%��-��J�^����w�!-'IB�h�ݣ*0!b�J\�ސ�׺�ŬV�{m�z�W��ށ(���r�R�+�'��
y�xR�[x\��?�I�ѻ�<8Z�qAs�;����/�;����f�ʮ�͎T��x�n4S�*S��Coԭ���������T�v͝E�#l��u_������{����
��l�"��}d7�*)��7�TոY�}�pԒ�a���BH�k�x&ƥLϱm$�b|Q�$+���{-�e��䯞]��4/|.������+^ԇ;�_ĄY3�H��o��.hC�Tl�&|k�+�d��_��������T����8��.����3��1���S���3c�⅞�`<z{��󗬗f� ��ڬƨh��\oT1�t���_��|�C	�w��_�L"V@{�hʐ��)`�\����4ՙm��|Cj�zix�5�X1��ܴe��8ҨU�����O�#�$�:��P����.��@���j�uO5�o'�n���Wa'W=)�����������mL��<f�9k=��
�\��d�ϘA�hJ�b�:�=lq��6[Y�P��~��[��?��rm�����b��j�yn�s���?�£����*-��6��4�(�23��'��rFD��~p/\�� ���x���?���!�u&ݏz��h\��ş�Hkǝ�˳����,�+�*�Њ�7J��Ϸ��K���y.{�O��y�L�k�+ɱd��A�%�\Zz�Q!���c�b䠕(�m��H��Yt�q�Y>�!}E��ȡ��E�[��~F<���ZjU�x�y܀�� �j'�� �z��N�/��Ņ��W��1���������ߌ�
)�;kaZZ��Ӥp��w���*�P�����-Ԫ_�q�ػ���a�1׎�	�
;�a+�N�M����_�v᪖!�k_:�����b�d_l�������~-G��1[@%X�H�wb�ev��w��	�#��d��V|JV"���%�T�0`��֫�!��QS��aw�������T���ACR?�w�UU����v��S!�"W�+�������F�^Ç1s�oj<֠��Y���j�+�/�x��B�U���	䩍�q�X��u )��[��I�ܙ��Ad#�q��Cz18����%gm�g�ZD�\�Z�p�/s�$(��͂�}oéU܆��ÿ:g�>x��M�8�~뻗�!O��z�>�SJM���1��q���G����C$	�6��ȗ�4��)�4Ȇ�3�i�O��TX��S�-C��`ݫKK�Jk�g��^3��z��������$9_L��an��	f%6��E��*9ܒ��&��O��m1Fvᢷx3�� �����⇺��3�d�w�NeM�S:�v�#����<��>�H��I�;�7wZ�&&V�S �0A|���c�R�)o����C�'��1�Nۨ���d�CejK�P0��k��la	I� `zH�Yw�ѓ�0d@�g�)U	y?냉C��&�+z��4�,�?�.��W}%[[L�zo)ՠWύ#�;��n�8O���2N?Q0������] �1���Z�"�;�e�G�p@u�����,ǁΤ��
���0d��f���UV��L�)%�PO�0W��������2ř=�H����/�`�W>�˖��x� 7Xj݆��.v���ΉY<�CQ*�R�E���5nF������6��0�6�$6m���(���S~^���tml��� ��HB9M�S���atO��ls��`3�=��_����N����{���(�0Hfك���ps8�������9`�6톿8�_�b��J:y��u�Յ}Н�2a��3�Wm=�AC���	�[e0�dȄ��]���,�:�[���	u꽻"���R�&����Zʹ!j�������m�8�
���� ��C]�#՘/x^:�M��*�ͨ
}���= >IBt�-���ې_d�qY�5L�=h��Ep�{4$���I�*�	�\��͐�e2�ͥ,�Boz����
k7I�S���� �h��渁.�����9���OTCH'��**�r%�p�n�{c�	���M?�˝
�N$Yz���w[I�ly{qI(w��+��̃�_�i�,�����
�`G��T��t���S�!�4ˬ7�8I��nn�%���'��#PhV�%[�.�]�N�zܴZZ����+:�zK�SU7�sV��3o�<]��ޑSļ��ʗ��!�7�[��Z��I'����mpN���1��K���H=B��%ڄ�h!C�eyq�����^$��(q|��e�yl�xJ\�/�M������!����Zar��
����n�6ͅ�fn]�Z��Ⱦ:�w����.�������o�5G4Lù�`H>�Gھ��$�3�u��������[CЖ�J���q��\�&	�j�)��q߷�7}���49/B���~�,d]�{v_�L�3S��s�D��c���kCE�;̒Z���ti�`+A7N��
F����^�0O��T��	Fd 4��|�`p!K�x*�=.�8Y���N6�ʼ�n�NS�ETֻ!���`�S���R����Z��	����Pߖ]u�@/�������!HH ^�*�?�Y,���߰�B|�`�X����s��Y�A��Ԡ��3�,E�����e[�0l�A�#�Bǐ��~�!�f0���N1z:a�)��������\��q~p1��q
|c��E++�t�g�N�y�*x��w��S�n���;�����&��?�ֻ��Б?��kg<س��[Hn��\N��P�p����P��Ύ2b8�0���!=��v��ͽ�q�E,���Ir7|R��5��]�Ϗ��J���<���H��ج�D{퉯ז��$��$���)u� &n�9�{�|U�߇ٷx`�)wR�M
�+�+`n��;�.b�^�X!��~�d����)l���������/l���됞�d#�����<S�y���' �d���>��`��]�˼�mwR�0��T��;�=� ֛���8 Q�����#E[��uQ1�Xc��etGjh�o��o4�@!���2W�T��A���&��f׼�^O���AQ�]�W�OzP�R�R����t�C�[+��3U�b�ue��;r��PS�������M9t�X��,��D�SOK�:$�����N.Ů<t<�{{�w�T��"0 ������?�#���n�Ze�]�h��iL��A�o{}�6d�H�O�������o����|�lo��[aZN�h���z4x����H�Ε?��}��!d�%�L�.����vT����s���ѹLh����xP(��u�:	KUKq�3�R�i����(���1���<�`i�� ��ɼq(�G�Ĕ5f�t<��O�6��R��G�`�l�Op|)�S\�}Z�-0�f��� 2x��xAr���~ K肏�9���1;>���V9 >w�G/v�1��<S�צDnq	Y%��e� [�($�႟��?ʛɶ@,�6�fCk �dF3�ve�/G�z����0FxA���
�M,Τ�A��K@*~|O��=?��ԘѼ������|�[S�AT���1�SY[{N����^W镖\Ù|E12����A��q��d�X�Y��Oݷ��I2�Ӝ�;w���}���܊	���.��?��7��m=6���#MU�hN,ȁvy<y�u ��$;������΅����k��9J5y��M.t�Z޻�ؐ�s����8~�=�Đ���4x?C�:m[(a�Qq�kEt�'إ�-�H��j��ׁ���*����*iW�f��җ��!]ˠ��"�}��}$0�m��L������>���(8���Jǟj���48�5�5��[���mAy��P�}����ǜ�񖮺���ȇE��rG�}�����^����S�GJ_ik���*�;}�|��Ч\z�<�ĝ�رAȱ2�W�������w��o��_E�zI������i�lۉ@-zx{_:�"�.�*�M$aES[A��G0{v�.��/�����z�q%77�A3��y�F�l�{O	��h�ak���u���Tw��VÑ���ka$�r����J&f�[tØ�^r���fQJ��L��"z����A��F��p��N*����~,�FH]�� V�1��)8�赃ƾ�Gq�D����U;��Q�M"�����n�֮-�0��$�A�K'�҇�x ���w�����<)u5�_�lKj�T��2�'���Žd�`C����F�_��BQ�Eۼ��̽��t�ox���:�zve�d�^�`��e�9�yA���7����9�4�o8��R.{�G7��al��=��勽AJ;�ɮzˏ��=(2��C[n��u3���.&��Y��N��n����Vf{���=�Ho_��d����,!�&�L{}-���7%m��!�e���=��� c�w�f����?XB��a���q�F �l�.��k�M��G;������{���!�B����)�Y�X[���jF2�谙�}˸��Z�\S������a1�I틅�d����)��x�R�R�3��cL�6R/KlU�)}�@G۹��j-ҥ�n�_�WiU�7��.��a`��i���A����"��`0=����5�ʖm��57��"���7�ӓ���ԶY��',y��L,C5+�˝�Ú,be�0�
~ᢸ�+J���Kyjmbw�d�c=Q���bw��=e|	e	e���eF�O␋�N.b���e�m�F�/U�گ��x{%D ��U�ʍ���p���Μ�r��s)(ҀX,żfm�p�5��p�[�$k��'4T�jl���Ӻbt7����OkEΔ�j�����E�7l�[��;�|d����A�(<t�
e��/�@�i�x�T�6�-��?�(���Lr]�� �恝j��ҋJǥ�5�sm���X~�	�/�`g�����:Z��uI�9{7NܞbJ��kz�Zg��%C���'y	� ��j�j�Q뼴���1@B����x�y[6l@� �M�?�r��<˄�J6#i���O��rX�s��o�q�F���D���~�f"�������rs��$����l���#�Jzb@�C��³dlZ�H���g��'�+݃��� �1D�>�ɨ�Ve��Q��d5�٨�;{%��~���=�����m��,Y��rb�s�)���s�������X� D�YCŊ Sd�9�E*��j��A��-�N�u8<: C�
�:��\�3~�R�\�w�X4�E���Ua�5y%n��Dy�ǟ�hiZ,����g������C�α����8��>xD�汢��r�㰡�x��È7�a_D�����N�jC�Ҩ�g@�a��x��pC-��^�I��|�W���0vD��DOX�:�^ �;�^b�6|���Ս5�4îAE�РǸ[�oR"g|ޔ�ޡ-A ���V��N(6t�+��?���\�L�= MjሺĆy,ĿȎ׬��H�dF?�?	x�Xe
G#nѝ2�Ll{����3����>���z�*����]6��S���3�^}��EN�5�,�bu����>%��Q���)2�j,���?����K��j�R�O	@L8�*��v�˥t�*!V8%���ᢳ�.
�e�a�r#��U�N9�T�?`ё��A^(�TNO��G����g�;�ê�\�� �9�$q,;�#���~^�u@�4�}��E�%�l%R�N���~�l���S�X�TACIR��w���H���TC�O��"w�t��lP\M(�C�*P�>��В��<{��n#� �7�M�5χuFY3�U������B��²ޖC5�͓����=Z�8{n�83id:D�%����^N��C��4��z�� U�o��X�;u��KFX\�F:���@�r��טfB�}&pB$�|��g4�Fb�PqV���>��u����'��6�ś�F�������F,�~.�eF�hh�$��b�p���LO��߼�6�g�v{����9k�*�h��P�YK����E�.\�nȦ�O�Tx�~lI^C�fwA��آ����ù2H/� kMߚ��;G��|B_�VO���^�Ng@�q�~�:�A��Ԑ^X� �TV���5�涣�{7��:omZ�;�$�x)]7Z�I&��� ���_��u��>� �Nד��Խ�7�����#@K��g\�[�g���{����N��1	��UcB��c� 	�.���8i Mm�A|N�\�cm���OǦ�x�M�~�U�I?�#�FzX��-d��"~!na�t9��u�$��`yL�;z�E�^�W�"p�c{�`z��8Cɍ��x
9���N�r�3y(Q�$��}k��UV`|$<g�O@�5S�Q~Z
R<��?��͌��NN��3hj�F��J�fG��0(x�\���o&1f�G��kq�_��Ԩ�c��)I,Q'��l4Ϣ�'8F\�S��x�Y��ց�%5:�5q��D%T�_��2��2�m�,7�eTv��PlF��u����;��N��)!�e���i�,�9��fV��xZ���]����q+��Vֆ=����=���,k$���ϣg_��R��bO)�v�7?�Cew����
�=�3�>�_w��J��$�b��^�c������(��qTՊ�x��,v�j� ��p'�����,��L���Gz�UM;�P$�1?>1����Y�1�\�����B�M9 _ �z�qc�]�o���P5#Ɉx��q������ϸ$r��I:�n�K�� � �'���|cٛ1��M�h
]�BOxL�e���cM����k��7�#8H��bc�&��~>s�X�M[I:��x��Щ|	"�����b�Em�F\s�X�c�Zg>� � @o��dђ�#�c��A$�h%vp<fBjG�_�^oy���`�6�
x�Y_x�����/�x'��S�{0�kr�Q<v�	rGz�(�U߼��a�X��h?�]X�1�xL�egw\�H?@M�0ܥ���
d��m�K�/�"C��s��?�&���}_�^����%;�#�AW��kщ��O��ϵvT>��f�Mhw��=�`9��j4� �f�q��θ"R���[�c����ɍp�K�@� �4,c��>T`�w�y|���6�O�+�)=8�y�~�{y#�$@r��g�k�:� �Ha�	ĊShѤe|s4�O<��&s<���d�a���b����d/��t	� ��D��WF����<����&�!���q�قd d� �%�UH�S��-~9ʧc���S'AͥݤZ㌲`M`d��b�c!e�K�؎m�2:�*<�w��00���~IpH��_�h����*���(�W��sg���JۦO_��݇�x'4G:�Eg���#LԮW��D�"j����Բ�0{Ҍ�Y(\5"(��ϭs�HE�d�]�{��H���ܾ��cZ�o{����¦6�� �r:	��Pt2B�?���BG0ߨ��L�>�+����N�J,S�P���wi�w~���3p_�������ѡ�(t/W�8��Y�����Ь֘kؑ3#]�u�՘����}�̶loc?OR���C�G�O�G�qܯ��jJP��u�Weҫ�d�[�8�;��\&��
3�
)��H��vh�rh!unC.�}��H�J�`�,�o�7s�g/��($��R��ݙtM�{|�UȰ��;>�G@���zȞg�R9N�3�LsӚ���O'ْ|��:��pU�!WQ�c�͇���&��R� f&��煱w!�c�k�NE���[�dJ;�D��)y�=��b���yl�.�#�<tαή�UH^9�x#.,��bL�J�0J`Ш|��5�g��E�"��[��SY����O����O�c����Ɂ��ҥ�V!�rHX��#�D'#,^�8<!1�\K*�Cl�L�\�?�����'��g���ۣv	>�9����\��s��hѸ&v\�^<�E����i�ܞ�ܭ�=�,K�NŻ	ՍM�
X�2��c����T{��o�'�Y��@G��)�dٽ�3Jl��7�o~\l'Z�tg!�u�:�˖p�o��6�(o��#�/�b$�o�a�����}�C�!Ǳ�
�~z.���"_�e���L�d�LS��vN1�iYbe�:���B�ېM5��l'��C^�t`��R#���c7ǚ�	R�.[\U\-�A��n�Eq�R��Z\�!D��u�q�G�I:���H�%��0�x�v���tx�	��p���'���i��8I�.�}�����;�ة��ԇI��cB��L 悎�u���=��*l�u���k"��r,�Fg�ld��_�##k�n���[4;
<>�O�LOG����O�Ȭ�����-[S�՞�:�Ѭ�ֆ�:n��#e��>Z�4�f����W�����a`-�6I�#9�C��c0��e�W��M�c��:�6�bk��}������u		,��yT!�g�Ƹ��9-�`�\�����k���A��F���>>�1)f���o���x�o�_��C��p�ݒ�X���-N���u񙼺���}O�r�N�Th��$:d�՚J�yJ�=�� �h�x�6V�/�H�B9`�qƏ�eϚ�������)F5�P*z��+��ڬ�Z����	���W}�l��y\�F�=J�������$:^�*df��fP�Pv��`�@D�#�S^MMs��>�G1���B/\���=�sPf��2~keĮQڤ�����C�~:�<�	�Bۀ$�����q�5Hux��fD���u�-?�DD7��a�5Θ��L�D��ko��Z��kӹc�rpuE�"�*�L����,b�`V�vۤ�"p�7��>�}��*�j�-v6���̍�N�c�9�Ӱ�
�o��&�!���t����M��9$�=�JL���U�0r��f�/�B��S�:1 i:���x�'�U-��@m�j�D
¡�LOkw�7jO��Ҷ��5U��-�|�B@��Cջ�YX6Ƀ^�t�m��=,rЈ�5"8B�D���̈́&7��pA���2t¾w�����q�	Io����0� �e���p����gz۳"��5��Lr�\�O��d抺άm���K�n�����Gm�.����N@���8���z�Sxl�=���:q* |2]�#&�_0�@�?n v�"j�K~w��e択נ8�B�+5���V��&	� �[$Ls�j�x69醤N�-��d��2��3�o�-�\8J��� �Ya�΀(X�F�-�g����	h�6���c�eF;�ִV𹌺<+۬��K���P�j(�F�����]����F�� ����Q����R]�+(щ��5�e}k��}�ˠ��V�M�|=	��Z�/.���!�A� 0�>��X4�P<�*j�Y������8�)���܅���m�7���27�V0�GȐ�,}+|h4��x[{�#;.O�H �d"�F/9��f=�e����[��d���(6݈��n�L��l�Ѯ�`�ܢ3���˳��dʇ��m�C�?�܁�8�qH�Q�r�u���q����Q�i)�M-�����1j�*5�K� ��f*�Ү7�5�IԨ������:���k�JdU���;��=?-Y�4˻�3�B'�.w�9;��5A��S�+7}��ۍXs�����TD<`7`�\\ľhu/�7�B�G�b�_o\mXl5!-y����u�֒��V�,�� ������P�y�($Y�"/��{���U˫id�
��ic�QD��,�lW��xß;�+6$S�dנج��|��D����Xn�������"��Z= ��r�ѨVn��5M1��[<�G��^���:�/Q�<�-g�����_�=�طf�D0q��E��vmmb[|�_���E.�#�T�>=6��)>�9���\�ڕ�K���[/����<M��`�qs�Y�#�s�I���Ii��b���6*�N\b��E�Ȣꤴ̡	'Bz-Q��@�F��+������
'g���V��>uJ��J�����!L6��˞���sV��ͳ��=��q@r��4��Nv�q���,�옓��)��ڤ{�UXA!��:�̢o)6�Cbof7v�!Z2\�&E*��y����^{Ѕ�i�@= tv�P�T�)}N�`�:e��X�+��ۡ$�p�FՉ#��(8���3�s�w"b�K�n�3�u�]����!﫳���L�A��E+�ף�ﴙ6#���0��x�O�9�U_f���sU��x����l�N�)UP�2Y�v���\��𰈷������=M�c��ob��<�P+��!h�=��������3�LR�w��Y�w٬��O����ElD���W��%1w=�xx2]J��O�`�l'u����e���z^SJ���uV�=-+�f�D��M�X�]���n�K�,"�>Y����e7g�P�l�;�]�7��O�h��HÀT�E,��!i ���h%���%��L�B�Ÿ�J���C�"�AÞ���~'l�&ʩ�H `��Hx�Q$�\m/�dR����i���d�}%Y?�t��~5�;�S��m�h^��R��W!��	l�Kٛ�F���� ��� ��1Qu4��}m�ȿ-ߤu$�CZˏ��!�˞i��~���b�vU�+R�_��i
_�	*Ǩ�_��V���+՞x�H�$;�98�,]�u�6J�.�����8jz򠢰����b����%?O3��@�i���y��9�#������m�(P�)93�gG�)0�"浮��J����7��L�6�A W�)�.ڿq��Z��d<J�����z"Z��k�_��i4�\c�F�&��'�>̷�j��rޫ���9%�?�&Q�*=�0�<G�	���d|
̷y�]��*�ua���oy�RQ��F��$u+����!G?���댉,`0��� ��h�]`�,��a)����������q^����<��-�sʫ�=��U1O�����h�d�ǡ�TnRR1ߐ�J);T�05�c�[@�n�.-i|T�>|elX�t��w�R
"�>mzʇ�j��r�d3��3�oƟ��	�Y7C��$�����]����L��ɴ1'�g��S�R|�sF�ܓ}�V����)�פa�V�P�'��U�C�(q� ֱ���r��n���r�n��o��0�N�C���$��v�`"\��-�4���}�7��t�>��v{���+3��?pW�Uc5�pˬ,dc�otC��#6��n�K�԰���ph��Do���"��eOɞ0�ho���aB̰����v�2J��ܞ圇�Ey�z��ݹR�����-��E{�"�CK("��p�f��4�2�����}���C�ЙD�Z���{��.Qc���@Ǐ��qϲ�n����a��	��V�{���]=�#�L ����B7�kZ�L �Ȥ�#�<�+��T�	 B����543��Ē'���6PD<͉o�^��=�|b��g���|ɏ�;�j���[t�rRoa�Ȧ���� A9���u9�Bc(�@(�h�6�/�ȧR�G	"�[=��u����\�Cz�/�>���!����Z�`U��r@���'�*
 f5��>���ȁ,���._�|`��%��W�8a��ދ�j5Ef�x�-��5
�����["��M�&@�!ǔ��_R�x.��@�lGo���������U�ҕ@�.�8&�S��QA�Z=%:��	T���w�E`�or�Lv��.",�V�\��w��q���<� �c%�ӭՔ�M�Pm?�a�@��udT�j�vl�����
���7��I\�����pJ�`���m�]��D���7�a��u�qH�"O;��hY�k�MѢ�
�<�)8>Bxo���s_%�l[<����Z�Ŷ1?oJ[��MT�݊�	�f�4�0&Jz���C��%O�7B�FY���M�4>']�)�'�#�T�C%�`t4_s�ր�kH_;=��0�e�gX�x�=�|�Ѓ�$��/c���P�)/���~-rZ}��B���c���b癓T�<nj�#39%?�Q^;E���NYF��K�c�A�/��q9bĉ�끄�GH�E1���1a �yN�D�*��ީ����y��}���
��Tl
V:���6�q�yCr�(^�?+F�K��k7d�z	�Θ�!`��W3��qFE�'
s�o�(�n�HOv
M�c*�zћ�-���.�UC��{�RG rA5R���3�X�����!hå�c~#�{O���L�cK�����C`-���ք[1UVT�/;��֝��_Iȭ��o�<9K�_J�дQ����������i��l7��St��N
qQ%�͡D ���.���Y��u{�p�@9ud�Z�l��*�1e	a��u���N�f%�����>��X86Xa`���X=߷��A��8�n�����p�5�F���K�z�roy��8_�D[�$���������-t�94�����q�ش2�P`�D >�Ǽ�1Ɉ��D2��ږ�A��꧅�rn�����b�6b�q��8��U��}\\09��E,���C!��:v� �2U!
Pxغ��d���ž�;���7�QM�@$���s|�j�4�|�d�-x���5�v��?oo�A+��Q�n�+9ص���00�`5�;�zيV4u�Ti�x�A�[� ���+ �uP��g��Q���9���	Zw��c�:�&�u�(��Sa�t�h!���-s���\^l�7����O���n�Ǘ���c������D4�<N󒔱��k�Cxdÿ e���0�M!���MPwŀ���a_�zvm<����b	t' U�!:�t�X�{~Ř&�a��R9q�:,��gGۨk;ٜ!�5-rY��W
��O|n9Ғц�iP����)e�CU�F��`���8�a[��;b�2�dg��r���aj*������>�e��x��G$.4���\�Y#v��f��yg7J1��-C]x��U�گ�9R_.���&5��PPIL��EB�:,`����^����;�=��{�y`|x��r�&�m�CD�]0r�ںX�~:�RC�K�Fn]����k��Xc���UX&�s��4�Q����Wc6����
��,�v���zj�(he!:jپg����,f�Eh�wPV�+��ń�����'Ws�\������Lr�vu�zԗ���AQ#K�=��P����+z=FOW�.�!��gY)�b�4����	 �+&�m�E����� H�W�I�AY�eVg�\�d�vMm��p��s	)����m�;k���Y�*��B���@}WD���}�u:��ɳ]�l���-���M6�k�ln�u(��+9	^��2X��uEq�xVN�]�7�eA�j�O�`'�,&H���=p6d���[C)[>��XY	��6�Yޛ& +Y�$a(���4������o~KF�@�S�[���@Y�Z����'��ZH�%�S�l���э�����=F'˘�P9E�j᥵�.#j����\��g����9�܇,E,Z�wM�{�ϱ��@%n�w��r�' as�[0����w��7e&�6�/zk��߲�Av�!��t�)���}�Sf�ܦ��*ԄN�Zwb_4�?=f'c���yhw�����D(T^e�	�ik�ki)�֝�%z� �\�+_�3U�2sʧF�A�b����إM��'A{?��rǜ���Y����Է�"w�����q�ѷ1���فn(��%��DV��4m��xf
Mi��b��Y�$!� ���c�ԟ�rM�Wɨ�C'0��Gh?(3fe��&Ҽj�dEm����M�/��dX���}&�f���Fۦ�#'��g^�.]�L�c�?̫��D�47��!�B��:�3�*ZC��v����$� 3������H�b:�����8\u02jK�����!�#jK;�<�*y��Ԧ`P�Y��'a�9Ը��%�^[�-�"��	�v�=3�k��D�pJ� ��b��l5�h�bpwx���e�ޏ�=?����������4�ɭ#�ZW���"��9�Tb%��TXf�Vk>�wA�5�QB�c�����2�-U�$m���mW~��R�BA
񽷠ɹ74_���=?���Z�'��@����č�(OW�����H�n<�i�Z��ד��-�P��#m6	�+s�ԃ�{��1G�����P5�mH���\|��F�ꮙ�ߋ�2�>F9�&pC�j����2�l����6��N����=����%�O�zT�>�b�ʧ}k� ��,��O��Ŧ�[�P	D��L�����b$�˽G���d%���k)��H�^��:>S�K�2����乵ņ�ݣ�.aE+;�
�3�8{��KR���x~��:5�*I^"��
yvTE��]ѯ��V5,�д,9��L�bH{g��=�U:e�y�q�@�D��ߒ�������Q4eS�,]N X+��C�c{{�D�8&�k���(���/!�,���yqM'�n�Dr��e(�Mv�'����Lu�'u�j��+Vh��2Yh݄�'�s�3�Ar�[q ҧl*<��9~զ���dM(kfqY��Q��84}���.L'{߽�7��)���+�P�k�dW������6�rJsS�6y���:;���U�3#�5���܋�3PΓ�����7�v��\�מ����q�����x��>�c�9��� �W��� 6K^��a�g�z��9if�u^dt�B����J�f
Bza���̂/d�y,���c(�����S��1V�.)��`n�q��8k{�6������GK��*��/�ɞ+^�s��q��Ь]%Io��,Gt9�e���m�>ބ{�n��ؓ#}Wsz���" ߞJ������;���=�A��rAy2L	�����-�+vE�6@���b�K�r���MDJ2M��2\c� �^���������Z�<�
~,��kC;So|b����g,���?pp:��}Qu���8�S�Z%�$$$�S�����(g�jQ����@"�3P��#L�&�9��p�I�V��,0��L`�	9;�S
ňm��~P�w��i��D>��K�E��G���>26�˾W���Vz{��B�W���TpV$��{��6
v>Ag��h�=6m�\��#���;���k��\�1ЗO��K@[�0��,B����t������@�Fx,Ԟb�Ԡ6�)=���Q'LA$;��̪{0��7�ʏ8�1uSN >�:A�&݁����H�UHs.���SQ�h��,�_�d%���>��%���g��k*3V���8>� �듊�]�}W�����O}����t7c��<C�pUM�`�%����rZ�Y�js���B��U��3�����U_2!�����	���I�cS�9��|���`��&,(GfAb�t]��w	��y��/,6��0۱��ï2�Xj<,�����ydB�T�?��V�\/F��]�2���@8�O�	��:閯�s�u���*���o6J�D��\'ךX��'>SrR�\�^��*_���&�a�� �5�rˉ�x�:�~��L�c-��a���V�vI��Y��$�Zїa��V~d2�9�>�&��[k�[y���u�;�i�T�&2����
��5���S0�d�@a^y���+'F6A���孚���m����7�X�\��������F�+����G���D8q���b�7m�ڊ&�^MBHԹ�+6��������4 W�_9r7z�cφ�VO�0�a�<��?X`[Ϡ�H�-f��ӈ�V�w���]I�>� c���B���r^�]�G� ��Ժr��d��� 9��9���_�ZEl�;�!Moc��x_S��������P���vvt����sm ��+2��3�Nȗ��J�?궓���)��Ig;,�z���� F|�L8�!J���4_��~T({o��zo��~d����}����vw�U�_���O_�VK��?A� ]��dx��!ui�C�%���j�CkCπ!�@Gh�?\tQ��c*i��;�).s%m��T|����Oӕw�u���Ǌ�,��H|C�{懳lJ���e�u	/�-�LH�}į
�^�*��ʫ��֐���ޅ]jv_+�­@��U��b�rx��g�v���p�ݺ��+�5x�����'݂fG0�`H������0�R����Q�6�鶴�6fR5��V��^WU��`lE:(Tr�>�V~��M���=�Z7q:����V���:@�����RN-5�Kn��{n��!GqG�w^�T���W���#&Gw���d8"2^��ǻZχ��9y)(��D�/��ď�*J���r�� ���K�{����j�dҷ��`��t%������_9��b�1(X�<���ι�d;ۅ��m��9�.�{T��8�T~�,-nu����b����2�lR�Z�Ȃ���;eP�=v�ar�9+�e8e�j��3�kٸ#�C�cέ�Ԑ�[)��4@�;�
�;�Ӱ��+4�iU� �L
�t�g�����/���)h�����簉�jB��4�jf͓&k����{�sVo㓓�S̡��G]���(B��C����TZk4">u�p�=-�yjc�`j8��|��n��5��w-Xf;ݜO����mGb�B�0nE���34B�n(,�9c @�R�V*�F(-l��$U)��`�}��Q;p��ԋ��y�-�;��9՜�=�Y��Yr �E��ϗ3E$襽X��E5��E�]`Ѳ��$��}��_7�`����^�쿡괭�[*��AZ�n����҇M=X /c8R�gOHյ�9�<��EN���+9��(���(fbK��R��
P�x���X	i�u����Vn�Q�O�_��W�v�a �N�PLϴ��
L�\�Z��ƯX��֦)s/yV@�Y,��`3rM+B�5�La\��+,�z9���F���ŀ��ڶ��h)��x�[���L�<�+�ﶬ遆��y��������^�#�G��p�͵p~��mm���|7�l��;km�*�Z�h/I��t��v�� G�٪��Nv�i�d)!�]���zIZc���m�^�%�O0�����'���Ka�w��@.?��c�yE�AI??��Ē�.T^�����.��5�AkfR��D� ���y�"�t�џ�Z���8:?r�=�n�Mש��q):,��&���Ҍ��/�fx�8ܘB7��Gk�A��ЖVa2�e����N>�;��j��%�qg�ګ�In`�#Bk��G�T38!ȡ�I��[����P243��$�a�T_���ʽn�6")F@�y�w8_R�K@����g赬%��Lb���{����KL�����΢�ΜI��^�S�m�T�^�_`3��vA����&�Cl����S�����D��_����/:GT���g�J�B�>��
����p`�h"��`�		¡���0�w݊o�I�=�HCg�F��x��Q5�J�]�]�:ݓ>�n�^�""	�,�H*Z��y�s�f�Y���}^����Ί7��(ܚ}#�j,�]uk��c"���N��p�F�/��Ӥ�Q�@�ub�H�����G"m���ڙhs�$ 7���MSa������T�J��W��8]���\C�'�k���[B��6#�&UXL��	��^���B՗ ֑3��$�28�]��+�d>F�2D��6\��P3LY܃dMa}�f��]7�k��ލW�1�;����� ���w�ö��X0VS���USJ-�yy��c�&�*N���Y[�dP�^�^�Vd��������*�~f��V�#Sf�/SM:|��p���c���h�k��.��wt�'f��<ZCAz�Y�W�Ɇb��ʾ�*�3�L�aX@�t�O��G5 ��� <|	�s቉������Ֆ8���3EǦ�H��.^hNv
�:�lr�][�K#&�2o��|�_��<��gs�%�ǌY� �S����-�y ń��Ǟ��r��D�"��1�Rh��2�.����P�O��euc$�RCO}�K���^А���h�D��, "{�ܧ"�a���g^a��%�`W�@8��J����?An��� �����?����������)�&��\wr����8�'�-ik��� qKinYs����K1gj��	��o>�Ww�<��p	 ͹�'1^�_���6_cى���:�7^&�7�������
���4�9��K�n
��6Y�Rv��.vG�@Y����ӡ밻o��U_ �t�<y8�� �h�45R� �k��뿣����3���^f/�"@y����RB��s��yb���ᎉ���B�=#�o���^H����8���^��xt�;J����>a�k��=��O�sO���x�)�)gw5k��@�BPN��װ�C]F��!�CI��zF����H)��:y��[�����<O�-��o���+�s��M��E7�%�1��!��A�P�\o��i��5�YkPm�ʻr�kƾ[�W5��{�]��)�j�"���a�b�,�.�q����9��߅fL�vt��8�����lg�.���w{�B c/�����s�S8XjN���3u8���}��;�)/�۳Zh��'fWf���[����3�i��jJ�ݻ�m A�8V#�؊�����0[G�p���{lʹ� ���})W}���n���C�8��8].g����$�鬤g�s�� gR�Q���oPP���Rv5���b�}�����ʮ�)&�ݦ�HTR��hN�>��S��d`dI�!�"�=���`���bt��s-��Y=	�F�<D��\��q9�0��Y��"sDB����c����B'&�V)41���ٌ����}��o}�pdc�����؊?�J�:�9�(���oe�A[]�����%7q�}!�8baaE�j��JZ@�����у���]�D����ީ��ߣ��~��U�$�"���Q�������_���<���`En��&\�ڿ�3���X�L"�������y�Ϩ�� j��7k}���7���p����n��k;O��^؉�>4��՘����7�o��cK
WB����>��B�P�D���W�#W���{��F��k~�3�"�!�΋���S���f��x�B>��R���ey�>���hT���_��^F�A�
���@�%�r_�:�J]�!2�E�\Tb5tj�ʅ���{o��?o�k�7�^���b��4�|�������<\3��d#����-���r�ou�����i{�T9�&�5�m]���:�xFv<��9���r�<�c;�����t.:J ��l#L��)��/x���H7b���12�eU�GN���9����u�gW�]^lp��J�{�iUˎ��dUB��UG+�|����ŜKk��A=�U�{.�R��;���J�;�\�n���m"}�H7��ݳ��N�!���WŮgjr�W�B�E�� C��(�V�)�^����or��ߐ�V#��A	Ծ�f��A�Out��!�N�#�ŤR�_�tFs6�=X�U�M��g��, ���Z�_k��$�b�_p���X�C��nGAi
Ї`�Ą��r��� ��>I	�C�%�l�g����'9Y��!V�/s�R������x:P1.�-������@�t�\��;�x+�.�Gd�ix�Z��\بtK#Mb�w�?n]�����Z��t�@��T��?)ZsfFt�s�-�;��/X(��4+�"�����DjL��bQyn�5.����(1s^ᐣc$��Fw�/�y��)�A�lh����[�T�`F{����M�IQ�%���km_��b|}��mn�����7�ʀ��_�c����r��F���L��9շ���~*���	�S'�v�����3��r���(�m1�骯�p��8���W���Fġ�X�H��C���٭��Qx �R�.�ݯQ�6���q��\�#2_w�3��_U���H{��u�rW?��s0�\��k�E#TÒ��.N������9�0�Ri湚=Zh�%a��xCܬy��f�د�����k�������F�.FNc�Z�Q���J� �T����3G>Y~�R�HB˿5g�J�x:����AJ�Bq�A��,��b��y�q�6��Ke�� 3���3�V5PZ/o��B�����{ن���*���^R�
��pN�v�D0������Mu-ym�"/B�ełg���a������X-UsNC�u<&i�ƀ��t��E�Ζ���� ���`>������|W�X}
I� 3��K.�͔�[��Ff�|�a�mxC�wL,)�Z��]}s@V����.�	���5]9_�)%}�Ы�1���רϐ��7�o��%7&<�LcN!��&���C�`�p/�[]��ĊS(�~+�QVR���d݈���C+�z��vKk�"K$v1M����3���kK��߅P7Кi<�!�(1�Xv�B'��.���v��9?C) %�_`R6����*)p�=4)�g��A����Y�XBLʪ�~���m��wUR��|�w�4�w�הHo�����"'�J�o��^a3p���ȵ��6��S����Z�����Wkrf���^��"g�*!�tI�i��J�����Ί):y���6o@1���:��s�}ܦ>����r�I���Lõ�H�3`�6i����:y̴c����nІ���o��[�����/7�b;���~��A�������Y\"�7�+<����!VF���ퟬ�+�YV�*�8e���TOG�M���#��I7�̃��}�l�?(�R��.G�PK��u����9#���R��GL:�y��xf��Hܸ�6$_�C��5�N�*�Q��ǉ)����Q�S����W�gF��L������h�o(@M(�W��'��ՠ�:T~f_�����[��Vܕ�Q2�L�4���?�e3���t&ɵ@��.5��*���p�Y�?n.��Q��RHf�N�'��(�����j��� H��u �cذ"�U��gF��Iphk{��z���>�{bާ;�Yo�3�"�� ,�ǣa�����1�rG_b'�M�,�`��T:�ෟ����!�n�E�W���QG%{�׽w��L��_�Iy�I&3����F�&՟�~A0��ܽnAp��]{���h�X���s(����7������~zv~<U>+�W��(����9?�*h�r<T�W��W��[�
��<j�h��1���[t�"��ո?^ҕ|��o\Z���c[v�ǔpv�
�e��0Q�^@�����wI�����B�4E���|���`H���dF?����3��Q��GI�y���1��u��)(a�ɯ��rb�W�k!1�0���Y�E|����:Z�Xڏl�R��x1~ȹ��ʁ�"����!o�3�POh�P�����~W+�ޡ�ɥiXv�w�g�5'��A�:��!���w��os���l��É{4I�����c�=HP
�����Z�`�D5��!d��_�8)ؽ�C��9��Cj��¬�M�˕��_��Y-�t����M�&��>��.��:�'pb��v�S9��zq4���b��n���!V�`�}ʥ1�8��VGb�)����vTk��N&=5� �aح�{����|��?��0{��Ő{����Ψ[���GG���T��P�n����L�m�J��rc�<��tG��W�_��2~�����ۿ;87�Q�;�)u�QCwnw\F��b�N8�&�P���*��Hd����I�{D}H��e�����~�2���p�E�0���0�.�㪴��_��xKZ����e�+G�}�\d�T�-��|r�J+���e�<�ZI׭ :�s~�a�v"��� tK��5E&�&	p���nx�4 ų��D�HlO�q�4F[3��`	+�Y�J:�,6��ꋭ���^�g��3cB��䏁�
T@���考cuǾ�Ӹq������T��J#1���C{��t��c��D쾈x��n7�Jj���L���p��/�n�n�Lm�I�z~�sb�;v��g��kX7�C���1��M�[l�}}K���x@!���xj���.$��lM�<��6 -��?D.12	�͎��8�x1�o��H����[p��tb/���m�@�bghL�Lkn�����s�L�P��H�7ir`Z�����t�e\���o��|����D�H�Be�+�+����H� ��K 0����&1�VwPc2g���j������S�k�H�	)+�LAYҕh
y@L����,D���ܠ/�M"|�'�6�"K]�����j@�q��Q�/b$��/�dq�	/�.x �匨��B����p� �~\x2�c��	�F�dq����1.��3��|v�"�ϻH[�4��7��& 1V$�/3�٢�v���p���r����k���ޡ'�@�=Z/�_�	<KjW?Wx�> ��air��١��;V�|��e�9�g�$Z.�+����	�n�D��%��?�;Z{�R4���?���x�T�񅽆����ޮ��,�Y^��FQ1)Z��6*[��8�e�ɑ��C��O��8j��x���H�1+�V9������cd'S|�<��	J��{V�x{���6���7l��]�=���3SE��n>?���9�Ml����^�"���V�󲶏]��U�?\t���o�9����Uo�t@��0���j�,�7�CY�Ⱦ3�q{3�]1j�	64<� �B/Ɩ�G�n�HHu3�F)��';��)9�J�VǾ�������kƋ�����i�kv�s��`M�E� bF�@�Ԣ�iAѼ�ݥ����A�����}��� �<�Ä�8��?
LR�:�R~�_�|"�)5�X��,\���5�I��b���6�3��v�7[T�ԍ;j��3~�{.��胿ӌ!�s.�`mLFH;-=�ָ�λG��(�s=X���:jj9��Hr����t[�%�>=u������.-�O>���}�t��2_A�ؼN"�����
Y�p̓��NA�t�sV��;���%�H���aj�x���g�.����׃�,H!ZQK��Ҷ�i�C�v8��B��f#���3b 5����*��6��yz�[��ME�ʛ֭�����gT����>������}��{V DZ��p�	�c��ࣼ:8�U�歝n*8��=��so'���/xo�{U�@T��[�jlaK��)8��ˆ5Yá�R��1#}Iyق <���R���h���O�?c�i�Ϣ�0/�e�,�z\N�>�g�xR���!6�<�Bf�	���cv1Y�ذ��lտKQ��T��#�!)c��.}�d�~y����K���?�a9�~Iu̐�+�ވ��"�i�=��~�ޓJ5v��J�,'�c"?#�"���L���.;b��!4��@�|ye �8m�P�<qcP�Cx: Ai�^�2��(1�>#���-Tu/�M�p�j��7��^�/A�G���xJR�.���|N�n�)Ӈ�rŰ��.�y��Y�u��`�>ϔu�M��0��_�p�-�J�{�8]j�����7{�U:��c]E�9cO�Wꄪ�6��w�؂1����lg�_u��]�xE.��B�s�`Y�JK"��n0T?:�{�_�1��u�Lml���l�K�����g:����j�AS�6"�:zY�ݞ��?�A�MW�*P�1i�p#~�
H�K֯��yֶQ��	���T�)戭al����8�q�'�����!8�:e�$c�X��m���_(�/�^���늳�;�"d�IZ���Ă�����F���BJfB��;m�,���?��{~\̹?oҗxˆ�k12"��H	7�,+��Ѽ��=��k�^�!���������Dkty`��ܸ�����`�rB|�	U��M� ��7Ov�+�[k�(�N���,˦����+M��#uM|��8��Z�h�J�X2W�t�(�f�V��5�,P�qh���]S1�ʎ�k�NI�;P���+��|���8�L��)�[�G$%�{!��O�����.�(fd���H�g��� >�,\� GV�ќ�gH��̡Jl1ET�>v	���Ox� FP�p��Z`��hR�ՎA�C��- �K[�!�H�S��Z�x���F�f�nS5�{�78/��H:��T����lgh.�a�2�c�9�UM��E���)���83�i���An��Ͼ�j�k����z�˛$���}�Vfܬ��$a��ߴ\���~i�B�	�F¡��J%6I"���H�t��Vh�4Ԫ|f&1"P ]�W����2�W��.w�,�a�܃�F�Gu��<�]�m���;�q��w��P$F���;1��\T�n�"��1>:�q}�N�p�J�?�c!�c����*���#2�/�ɒ�"N���	��GN�b���C�w�!p��U�ԛBXFX>�>K��I|�'jS���a;�s= ��E5�n�քE��,L2=+��lKu�$��7�v��9�ש�֞GG��T��wkPV/-y��_�m���������qP��g���逃p�>���b��T���#/GĦ�O:�^��	�
�}��"N��
��J�e��q���
1FYZO�)�u�ޔ���_}��zI��E���C�����A!����xjǞQH��cä1��(~��ux�B@%���l�/�C�V�(�P����� ���/�6�]��l����^���� Y��e���1�~#�*�E�l����wU))�i�aF��h��j�#�Ⅸ�idٙ�_���P%F�e���,����&R?nv������R���8�pp\h���jZ ��z�="�{5�P]<c9 s��
'�0hs:G0�kf���8�Hy���C�7eƯ�S�(J�%����r(�$~ϥŒv�t���]��͒"v��1�_/Xo4��΁����6e�5��~���dJ;�_:Un�� ���.gs�矨��;e��;�g��ך�X�����̷6�j�nk�U�"W�4���կ�z:���)uC��,���ϋiX�:�פ��G�J!pB����?�33k���R�!)�}�5�PZ�u�\E�&H���Rk��G�l��f����-:
��m�$,]p�C��e�sz�D*`-q�5� .�~�s��:!֦Q�>i[��|�\���ItU�[�I��D�Ԋ7A����@͒#���c������?���bʕ���h�3e�̓s��f��bD�5�0��E����$/ �e����7�ڃ9�%�f�2�5�I�as"V(��d%��J���4��K����ы<����%��w��WD-��B�&��A=F��e�Z���Ņp�	H�E�
����m���̼ifib����e��8��uADUc�9Nj��3q�a���c�S�����0�=�o N�%�FF�Ky�����P'����F���<<ko�������vjP��ꋧ͒��w��4xJ���h/��!aЋhSw�,/�4D��q���*�$ڋ�
�5���zV�KX`��Yi5�Zؗ��ˁk�{���I����(���O�d`��Vc���qнSU��R|�R�Q�a��a�wӦo�"ʚ�H��1Ҝ�������)#T�z�v����g#��Y2��~&��,*���Ⴋb@���-b!?cf�� '߄P�lI׾��^/G���d�'�	�����65 ��백���¶m!�������5J���*&�'�ݵ�W�$b) ���ف�2��:����'��(ZSd~t]��� �2.��?ǹ��Շ´Vq�$�Ɖc&�|�F�}��g�LШD�~*���`b��b��ϏxI(٧6��p`"�͔�z�N�zv�?����M ��<�W8��>-�G�{��jo�,iɶm�,�/�~�t	h��Mny}{n�K�f�����Q� o�I�|k,σ�h=����B�Y����;duώ�W&���������ۅ�m�pN1.r��w¿K���2v��,DU�v�""M��(�ʽ)��ͭ�u�O8i�N;Ĺ�Q��ۼ�x�N�V�AؤS�_x	}���&�z�W9�7v^�����Y�m&�Y�~d�ٿ�u~�y��qZ��=��7��w�"�FYI��A�!\����{φA��E��oڗ��ƞψgX�����]g�Zd��,_1���Zn�:��A؉u,�������~|�殄  ��si�dߍx�2��Efq�J�)��{B�M1�}�ׄ?���{4��}��'�=�������;��;���68�Ņ��uՍT����&e������ >Ab�lD�m���%��]&I�.'}V���S�M��;!���(������Iv�=|A';$-�	�AΒ;���d����A��~��E��T)G�/O�
䙕��%ȣ�3��mm�2��/2�`����k�U��.�[`��__ї�
!�x<���)���N^��&���Y=ޚ�2+'c"�jF��M����5�1k-ĩ�U��:y��A�#(�ᙣY[a����7���$�atC�&��>�'6��f��
����>
��y�����
t2O��a�ܚH��R�j9�	�Qd�;}��MB���q.&����p�;:�0n��:0����M�I��b��O$g�9�
 HWߴb7[��cA~��W`]"j���T9�����ip]=D���#^1����	M���go���h�I�̓"%?$�!�s�>��@�~0�_���=����I�R4� )��2p$n�Pf!�D�g`����FKQ�r��e�?t��N~b��Г�����Ym�O�	��˙h���@\��j�܁!�uL+;��� �������Z=���s3����X�5)o~�J*�t:W٧���
���e@���.�D���I�l*�	&=���ysx�h�����>�������C>Φ�)ȏ�-\�FCy��)PHusw�ddj�.����F���mĘ��fpJJqi�ZQ�bRC��$�.,� �u����:�I��w5��Ɂ��mҿ��u^7�q�F語��J���'���$�D%�ľ�n㶞� ��vvZ��]N󍀷y��Cd�U`�VI.�A�b�3��˅�Y�VgKqp����� `�w�)1�n� �2��D���y���4�i�??l@!�R=-�	���lQ�
� X�]���<\��Cm�Ñ�_u��5Ԇ��?�80���%R��S�i��᏾)%��5u	�$7�t�0`e�9��������=�oܞ�oBt����i&������<���w{!'W��S�����5?�>Q7u7j�^�[!���Kk����&�?[�l��g�׭\��iG�5��JP� ���)+O�M�O�m��&(��UlliU��9^u���Q��I3ē?y|��ŀ��ųV�5!蛥_��I��h���o56hO'��
�RyJ��a�n佭�'�c����64��Y8��lx��>�+�$s1�7�n��ǋ-ͺ<�#v{�����(RK��K#uь������$��i>ƃ��������͊n��y��E�"�gm����c{\נ�H���)�����#��B�M���萸��TGy�����n�a�������}��':�X��O�jE���R�i	j��ժD�$ ���	�ѫqZ��U���.���4���bV��g
��DЪm{���`�X &�?[�.U	{%m�a�H��V���4oĵ�?u�(
��|o��ј#��#��)��X���ULwGL>����� �NH���ܟe؏��';z~�؝�c^L´)#���ɜ))�&�yB*N��PD��(LG�P�f�kNDi�L�Cd<*~��Y�k�-b'�컷����2�  M��*�����O��~��nV�B$�J��تW3/C�5T4��i�q;�A�_�#���A;�+�YWS�	7d�@ٍ>?�H��ۓv��R�G����R
��㖻��
ֈ�W��%����]3��_{�y<�*��vEl��U;�gu��2b��G�1�f�"����'p>�����Cx'�G!�|b��i�S]T����?�ߍ��9�f��[^����*0���I��h?}>����K���Y"C7�4��d"������`��v>�ʯ�� ��[�ws����ϛ�/�qȶ�����Fi�&�܎ۈ��o���%�ǃ����m��6�񔜃̫�M��KQё��%Z��������C��R�{��뱈l���ؤ5��z���?��{���<ļ�	\�#�;@��A��k��'*F�T�L�g�hT��d2��b��ӹ�b��E_	N@�4��'��h�?���m/ �ƃ�Ve���	�Hg�)`��s���r��p=��h� ؘ�M�n�3�I����z�� ?|4���K�m��jY�� ͟j&����*�TH/��Q�-�k�@4���jB\H]�9\ꁂ�끡v��y��q��Fw/d�/����r"��Evw���t�K)�=7wdd�+%ѡ��Z���t�v7�Y��O�n*�=�IU��X�g������u�H�߀c�Ŝ��A��F���kS����r#Ԉ�d��Au3�c�^/Jk��E.@�AgvZz�,�\뚅-�?���2"V�&k�Ȱw7��8��f2����eX��C<qMTy��� 1��,�_�n�΄��S��k�����Ɨ��e�5�����Tg��M��@�QhQ���\JDh	�P:L�6�6O+�c��3��ZGX�'���]���P��WKQ9�K�ڱ���
�e���Lu�����#s2�{r;�5l÷X��ڈ2��	�����x��N�􄖔D##Qk�MԶ���J�?���q�.���1��r��Fr�<�r^��o;�p��3�r� q1*�����K)�
��&\AQ/g<b1�#�>6�#W�:���	�w'O���V8N�׉�G�*���I)�(v\[F���ֺ����}���ۍ�ŷ���y�r�smh�c�,���ضO9L*�ud��2�ь_-/N?�xK���ҰP���-�@�Z-���x�m:&��I��ӽz�'l��W�@Ղ_u�Z&��ӂ�3�kkJ��\�4��� �e�d?j�9��R�	��N��e�A<T�q�����7�H+�b�a����TMiI�BJ`�w�oP"��Q��ӥr�A��h��㑺�h�ݤ`�'��W���?+y�1�.���۟�2�ɚ��m\Xk��R�:�ьv�UO?4N�-,b��B���c^�q���e�e��07���%���f��h�=ŏ3�ѭ�>l|�����@'���?�2;e�kbM��G���Y�����|���Y�������� V%���Ǔ��rӤ꧹�X�Q*�.�_e����]:��N�i��(�A�a��#��Y��nE\����cG��7�|=$�jH�G}�ƺN6aV4;��Ex����Ԇ�T�o���e�ʿ6��x灻�g�Cu{�������h�`^���m��̍3�b�fU�,>|;A5*4]R+Ufdד��T�����?�dV��-P�m̆�b+T�x���:�-�z/����s�4o���H#��)j�N���`�=�0����>�j��Yoչ*�Z账o�ш��y�[h�}�K.=ż|T�%��=�w�,|��qJjH���T�{��H�ʹi�u�AEQTmؼED�A6؟t���+�@�O�@��J���M�⺅�rkC��C`��Q��Xk�渚la��+��ƙ>��X�e�\޲��=�I��uo�7��vR�[n; g�B
�	.�+�j�G��4�#��{Ƹ	�]��[�uO��{=!|�^Uu
_����H���<��.'���gVNbq�t�C$U=԰���oӇ
�/�w�i9`��M���E�]g���9\U����Է��yy~0��x1�b�RB�����?��`NjB���<�1o�P��j�Y���S����=g�6 �X�х4��K{����j�-�)��Y49��>m��1C��4!~!�k�U�躓b�E�U��`������7�dN`�0!'���(5��DlGą�7mD��Τ�ϡ[ؖ���iP�U�(|����Ĳ�d*N��=F<����HP� }@ڞT �ϭfW�xU$N���, �&8zSx�܉˥�IZr�l�t��Vy��R�=�fQB��qw|^��|�.�t3�
��X<m�T����\��~��#����a�e͌����1���ֿ�V��5�}
GQe8���j^�I�]c��Z�*6/���#�=Iq̡��`{"X2R�q��Ų�N��c##gsY_-���:��|(HBs��uA*�y�<�|ʘ��Y��;�J�5�=�3'�E�
������6��*R}j%�3���H�C�ᖸY��0ſl��4".y��X#_������<�B���M�(���Q�=\)N�Z:��WLV���1��Sw�g��G�{�oWܜ���\�\���������βr9�0�<U}��G�/�tc�>1L^9k�|�%��<X�p�Wܾo��A2�Ă��N�<�B4��B*#oB�٪�E3���r
ir�%s�����r�հ��x2���7�]$� Z���� z��iz@����n�7j�:v��N����_3s���go╆'��?6�8�ts(��_�A3�f�)n^�E�I�H4W�Ȼ-m�����F7�śs� [,+Z4S���7b�1i;�a�|��O�]UaYxRؘ�J��{a����oG�!]��ʸ�š[B�X����g3��)��U�(d��B�i&עô���[^�e)/��~x.���eh�NI�3d!a ��>B?4w]�^�d%�D�J�,��Lغ7)�.�����.� �|f*�C�>	w�Ol?�1�3�X��*�o�wE0�%#&S;��L؀�RۑeR��)Bs �������jG� ��*�m��Y8f�&�iI�d/��"�0���?w�XfҀ��h�3��	١�k�̉y��@�ɸ'��Ʀ�� �K���C^Ӵ� _W�J�L���͝�������4�I����qj-���E�d�������s�)�ӿKj�Q"s�T�u�̥�Jg���[���aD�&��h�'�Dr'�^Y��`�.��#�|R�6����o���s�d��	+�;�x�g�^B��#��5;wzε:���QR��kJ����0
�z�����(�h.g>:�]�%Ρ��I��a���ʛ��Z�\�{�?1+.W����Ɓ%g��QhQ��3W��Yo��q�֋M.���
޲�\��PDi�<�v1�MC�q Έ�l��Z_�=��w�J4.U�?4��{J�<H�h�W?���p�����t~�͔~�-�<c�\�_��1����������g�-PV��oY���r��苊t��d�o��� ؅E�;V_��"�q����(��4Aƾwcdg��������R\�u�oS.��c}[��E,g��K�Bz�8��5ͮ���+�n6�-Q|�U�N�*o�H�J� |?���Sf�@��.������3̜}Fv�@,~+�77�A���N�+ۜ���\X�x�YGӱ�݁��4��75®��K�m���!IV�˗zI�@�~ۍ9)�p���
�=���$���k=�]Y��t�4 (?�`v�+�c�?�%Ѕ��S;G�0-F��5\�������H��<r�C��$<H�p����/���+ax�5aQ�E���1���_�+y�
��Y�F��N�p� �gt�Ѥ2�[��^krj���г��r+�W(��j�tx��i���or����Z t��>4�	�E1{�"���V��K"��n�Zd�^5�N� GUă!��U:Uv8���ao�Q� �p'2C�%�S�8��-��3�I�7�Τ�=O�ˎFo�T:��OhU��X� mFy� �|&L�x,C��P�%�5��B�õ+��*֏����w6�E�Q�^�0P�i+j *R�p�#Z��j�����L����`�7��A�9#߽gs��U%s�
oΫuC�S��G-戠öڎ�cTL9�$���y�)Za4]����-:; x��?����u`hy|�!���vlD�9/I�7.f�7��|�C<�J�#�m!S�a=�||����h2G�S�9�uԗ�Sā�D��ې`륷��
�&q����o����i̺k��C�8�K�T�'�����_������Y%>ވxYD��{s�*��>�,j{��cɆRq*�O������~-�&���a�����Lƾ
����J��>�V������÷������T�(�it�SG{��uq2�E�ݰJ�&�R"��] Kv��2�vFx>)��m���Md
W?�'윗_������=|���g�E4ē��� ��[>ܰb�(�ی��F@�"�h1IH��Ӿ����r�#ى�?I4,�bA殣���N�����6H=\N�Gk����"WJ�O�i�	�a�V�&�M���F�����*����tU��A7����*�D�{���2��z��ty��ZM{�&dh5��K�I�B�T�Nj�J��D�~_�=70<7�-G�(Hy�X��g��O1.�����F��uĒG}/T������qr�=I�`��N���z8r����x=͚�}w���8�N��o3�����P����&�7�D7��@`�F��X~Y��H�q�YD�����Q�f/�5�e��[�]V���Jۣ��B���W[�~K��Q��MM*%x|Y}�2I�M�鹇$,�IJ�Mغ�O��3�O�Hש`#�u��.ō	[f���R��-��JIw۟²�_E�+�\��{xr�ݨb	cּͪTK�&�z�^"�f�d�b2�{ npy�b�{qO��"��z$݋��cV�P_�=B����RB�Ffb�_����\�G3$s`K��*p�o/���72�����T��rB1���Ж�H�/��<��tǷw	5�"*���n�>��?Evҧ��qN�ċ{�����}�dʄ釧z�Tμ�OM&))���GM\���Ѧ�Ql�-�V���h�7�LG�6���������n/C����i�y،X�[���d��]�3��.��>�(TC[i��VU>��#l��`��R2U�}Ϡ���o����}WnRg~�K9x�}i��G�~���C4�Q�����Z������d�_�Y�ч���k ��������*�:�ǒSi����<D�LE���f6�@ ���FP~ۜj�Wz^}n�s;��{��@U�Ta�3��E��Ѝ�G�|m\���~�gP��J*f:g����#�m�ϭ�+e~����Iq�S.qn�Y.!Ml�J���+ʄ��;kt�ExH�1n�^܏\3us�r���]5C/$*�q�3��7	�]�����FP�m���9��"rpm���@�N�P����������qŗ�S��6��D�_D��o����BS�ז�匳oWoÿ
��f��[>i�Y� B��OI(L��zE���55g\O�$��c�#���n�eh!�p#�I��Q+
���̿f�
����	(Ғ8���F9��_�$�3#S�~��L��Sk��{�8�:K-��0@s���o�h�)f�(�:`GZ�y��+���9���`@�k��vլ�)�Z7��g+�׮�(�u��
����N
D�[���XU�����=��`�����6e��1���k�+:,K*TIv2��B����@ 8�Y���s�-Ǯ���N�M'&���^-+6�qAƧ�;����`�6%��;k�$���Y�p�c=�ϫL��D���/�?��|ܾ�A�n�.]�?�%�%B��6�5��)�J�N�l�v=Kx�xM(�<L!�C����#R`SJ	�)�
�`�����0+L|��} WQ�O7�cq�PmS*�r}xF�u~/��&��?�q���%�^�����!�I���>�w� ;&��z���.��~�������ό��'(�<c�U/�j� �M�*�p5��m0�T��1C����X�
��`�2�h!^N��a�7qnS&	��7p���T6?�N.�8 ��&b���r�b,�?��H��n޺* +H����f̦�^ƅ�/��X)�<����9�Wl�}�9�~�����\�(2G�$w+lZ�H��ފ9~��{K��z�d��jA?��ѲwgF�.��4q�VW��#�BX|�0�8rA�_���[[	�8U��`W~��XK�s�`z��\�Y��]|��n��qz�\�=��F%�`�4��BG�U�0]�dv���e-�83ݴ�����}�'�OU�������i���Nʥ%�g�7�Y�:+s�a5���i��t�Ճ+��Xh�_��!�x��v|���B�!�U2��P� 2���N[�m�.Y�D8Ĺڷ�f����DD�}�\�#��EG8+��Nv�}�"�cN��UIY0�շsp�EZ��7f4<?�2,aC��^
 Wβ8\l�C
%���vzq}�����?WC_��l�	�ט�_������1��w���:�Z��V��	sw����}��)5VT����>9�x�j��LH�k%�`Q�o�d�mv��B�asʱ��p���`Fڛ�H�o�II��*v��Hc���3�N�	T(�;��������Y�z���{�&Ne�k��DJ2/`�ۧ����W�-ae@(%7�u�\��:�|�~y���;��X�3��b���/��91q��u@�nu�v�d.����ْ�F
#�Y{~e<�a�Dގ���6��Z]-�ݲ�&�T�]�e�Z��D������K��^-y2�����F�m���TIԾ뀝Po�����@BD��vŠe�Ԭ��N�>D[q&u�6�o���`^-�?����m[A^�Y�d[����i���S�e�����/��M\���NB�vŷ�1�F�X/ʫ8�+Ԃ)�e�����[v*;>�k��S���UF�B
j�&y��~�R$�N�K �����J�^�S��1W�:�:��AT4��{ˣ��������X��:�k=��
��!�s��$w}u'ND�����oI�t��a�Qk���:��:*��}��L	n�b�S�����@ �cH��+B1�y�ǆ)�;�,���}��֔_���K��߰zO���.q)9��[�A�ؔ!M�G\���3��7��|c�)NF+`w�M�%��]�	��,Z���Cc�Ej�� O���և���Ae��u��
�RGqRT���&m��U�W���M(��m�V��Q���z'g֗Z2��K0�Yb�6��Yo�~˔�J%N�&�;����'�@�^�����HL��/�I�}�8�BDXK�13��T�c�������$^ ��v��l�c���i����	!�����������ނ���-o%����|A��D�3
���L'7��yJsUD���Dnӕ�C�n�<5R��bFi��c��w�29��K0C���Ș�.�dES��dH%r\늴�Q�>� =��m9m����F�W�M��<}� ��E`$���<����B�3	�۳ob8�[u�G����y�yv�ny�s]'�6�My�|բ1�r��U��"�4?����a.b�U4�#�{��2Ԍ��N�Y/���?���*"?�m���;�ͨ8[|_��5����P���������q:+|X�7"���ڴ*b�"���D�K���������%���M�h&������\�E� Y�Vt�Z�ՁK ���d��v�z�0����uW<$���#t���z��$,�`[��gF˗�$:X���B~zD&��=�]=��(sc$K�BX��T2�UG�Dʉ�?;����'|��H�wy}�����J��^�EX+��������m:��tͫ�����g�m{���V���V�N|0����s�K�xt�ѱvvg�#b*c�'�>(d�NE�F�9v0�����^�����d����ux1����6-�c�w�cy���L1�U���q���岙C8�}jIW��Ѭ$PtdG^]`�?eR;�*����J�����a��=<rU
Y�O�� U ��}`�o{��(�T� �b�Cbǫ\�D*tsn���������uu�$��>��<Xl��DR��,�Z(���I-^�c���N֝m���I��׏��MDBl���g�*A�E�9�
�U*��� .�g	
R��!@k��U�Ϭɛk��O���v��wFmf_��OHG����f��X��]��
u����tV2��BP��.����,3�pm��$N��j��e@��߭��zC���U�w�%�k����c������a<��h���7�B��Vs2����ֺ&B�y�yyr�J}��şJ�ZxN���h��.�����g�+�x���*���X����l�E�l�Q���d��5��B|�$��
�lb��%�ѯvzɐ��%)�i��ԟN��r[Nm��cH�|��i�49����y�u�-!ۊ	{@m�����=1�}X]���}��9	���)��;H��O����vƮa�X�=����?'��I�}gR��C|�Gt���[��|#���i	;#v�7����]��i�w!���ʌf�M�W4PK�a�{�v�=��xin��n0Lfq�9�2�ܾ�Ƹ�ו�u���4j͡.e8���A��a��A'���N��΅63Z�a%D[.���	I�Q���8T Se��I�(��M8��	<a�[jꩤ4�K"t�����z�ڡ`&���Zr�P
H��#>9�j����Dt�>�<��X_1�8h��&����Eo�h�����>�
��[���@B��Q��Bz�,�����JA��]���:J&JH�ų]K��B^�֫EO�5�t児��K��[X�mE:��)�ƛ��ЦSm��!(�(k�x���� �����b{��j��@��I:��V�6.��ў��o����Ɇ�^��@��	g��I�]�k+����0��ۋ.�r��׳�L1[�9����Գ�� �JKe&B��*���є���Wk_�,��YY�� �4��`��z�a(��j�N��*�������gȚ�]F�����b}MÎ�k���vl�k����N�h`���{p�Q�#	�@��ragc|�]\�l���%���
-:*���;xRZw��{<)�#�6�V�@/^�S�2%�� 2rM�O킛>1�93t�>�a��7���������W��-��g�c���c�RM�@�%��ف�J��U��/���������Om����5�t�Z���Gj�s�c�l�حݶ�D��z�C�������M+�R��*�����rl����w���NE9� _�r2�w�]��/ ��c���C����bHB��ˑ�%EwZ�P8� ^�%�t6_�%�\$4O�f���}�|�޿q��avB�����5&k�(ی.���#x�.��v����bꅵ�����GFٗ蛬��D��U����WF�쯗t�84�o� ��aS;"�_Y?g��:�C8T��r>��M̤qJM�a��荫�/}9��?"���@�T����v(ۑb�k�aY0��DR ��uȐ�t��3��+�ɃX+�ԢU	4���Ʉ"W]%gȪX�p1u�|�-l����L�pH��Nu�^M�+�_"ψ@�\�\���|���ْ��n,�l�J	?jL=�*�;��.ʕ�!ewJS� �\�fR^�6�P�����X��ʓ��n[�z���e�?I4��s��?�/وv^_{a��z�p��!9hLq�Qs hL�l?9q��(($T��g���ye�@�~�CR&hiZ�Wi���@�99Er�S��:r��T^KU�oE�Di�ך�穄��)��czql����՝�9UP��+J��JT�+��{�Y�IL �"���`��~�!���J�ٴ�Z}±���e���y&6v�4�q6m$�n������T�J{����~?�zlZـ����~+d���z5��=���^�Mr��S.]�{��#[�^��D��@�V�O�HՊ�:�q>t�]��ǎ�2|x�g-|�e�.�������rZQIh>�m{�h�2�zIE�kӗ'|�U��M^m.t�)i48�kQ��J�F�@�n�p�b�5���%u?\�IX� ��I-����E_���I� �j>,)Rt���"L_�+Ea3'm��v���mq���G#����E��-����zRǭ2�r����A7�R��#9B�c�)m�zj!2�����7&p���U��'BT�J*ɚ��$o8��<�Gx2�j���D57����*H���Mj�l�Z�������{Z��;Rڣ$*'ʌ+��$�B���:��T�����u�֠{E�~Uڈ��ũ� k�6b%��5����+�P�A�TU�y{�8Ηf��#�4��٤�^�jxYļ��j����ϱ�6Z��������Ӥs6�D!U�g�2�3��	����)��5�|��[λـ�
	\���k���ȽE�<�; �~�cG���*��A�t���[�I��2���b���[�!�QM��L�!��_�D�y���zݐ�����]쫒Ql�� �}e�z��7nC��s b=MF�CfD���2�mM��aD]=�e_<n�M�1���˕�ڶ�*�h�f��O$TL@\����XA�rO4��I.bQx����M)ff��,U�}Y �)_N\����{4�̇��Ɏ*FڇDڎf�ߏMx��ud�������wp�N9�#��c�J��3�?O�����q��g(����O6\�)���F�"x��dA�g_?�B�U#��K�d�����C�Ƚ=�9� z.n���;�Oc�����O��S�`�Rr:�+P;��T�jXu��Lq}���:�n7o��p��'�7��%G9I�t�0Q,I��Zb�`���6g�y��>|�y�؎�9���b�ܺ�񠯥T��S@`+�<�!2�q��Z�&67�g� ���ѳ慦#TF�e"����<#'�nB	8�Ca29tbVߣEŀ�ԌR��(,\�����6z4�Y��D��{�5����@޽���Z��l#T�:bafX�oX��墪|N����w]-�o^��x`�b�����5k�*�Re?�֊Y�GrO9I��Ђ0_�+x��DRսg@bE���&hD0�����247��ɸ����+�N�Ⱦ���W	�����E�n�Mk��Hd����5�m�4L�����N#:a���j�� �0l|NX&�?(q~�:�Ax?�P	��Ɵ��n�GV1���$�9.;l'��7�н�/���'H ��t��-Q����Ҏ�<�yd�6��g�����t��5A����͇�(��3�v3�M�����N
�rm�<�l��LQ��$�v���|�"��b4ذ��U�5���H���[i��wn.m"����Dĺ��c�QlV�v��}�!����ۣ�!��P����BT�k?;\u~/f��UV�+zE��S��8 ����21�?�E���H�P������@=	|rlI�z!k��|�:x�3ޔgI����[S���x^�LPq�u�̗y�G�?�}t��p"��8*#��ͦ5�Q�+��!���Ջd�����97xx~�����]�G������SdJ�[��+��y���Xv�پ��y��yP�* pj/�!����a�3O#bXh5�U��_�^r���^�!��̰E-j�:a���_뚒�7X2�{ޜԮ#3���
(qR[#��!�U�
��A��}�,_m�T_�s� �����!�	�z+D���b��m`mo�Y��"�Uf^F��ՋK� !��&.��5�3^rɼ�hy5��]�i�l;�����w8���S���i�4��O�.v��>u;���G�ER9a뛹WrY�e��V�;��b��a�`����x��"��zr`���%Zc��A����a�bqCX���?^!��s-A\b�p���Oc��D�=�!0���ꜨӖ�Sn@ï�;|jn�����U�N�kʐn.�W��g@u�E ����ޝ�F��Ӛ�*�G9�m�.(Ȝv[Q���4��L���19H}ճ���C�+0Zec��l9���#�ճ$���j�ܴn4�ys�L�Au�뻥O+���[��L�r��$'	
���%X*$yw�x<' �����Y�.'u4�����%Q�5�)����P*�z6�	�v`�N��ջ��
��`S��{��یի��q)uVcR�������fB��A�Um���1�:z�r��)v|.���0b��m֎`f&1||�/U��G����#�ƨ�$?P����0ϏKQ�V ��v���F�D�	��&��I��$ 3M���I%3�_鬲�]RA0p/�D���Ej�`�P�<	xX ����pD��,�.��Vu+�B�p��b|֌U4#NKcS�#]]�Ʋ�[gX���[�����5"�7�X�����N3xS׿{D
	^���>j���)�2A����J�JG�"6����B���]:�=���Sp����u4��G�C~��(��Ը�Om����)��f��[�Y��N�_��et��C�l�p�ݳ���i�������jLL�I�ڌ���(��	�O�AEy���d���IYl�Kܼ�U+SMcU�\j�'UQ��Ⱥ$���:�m�rS@�|�a�����n3֔���y�6��x�*���	,0|E�8�%+���Q�`��rt���Z;��v��QNK�ӎ�!R�L��zݱ*[@59��C\�Zfs�_F�?����?�곷�Y�^�S�(��o�I�|(�+�+
�tb^����pA��t�iBA���T䢟r�oaM>g8^��b?~��;ݶO$��ӡ�������Kj�gN�t!��pڸAԒ�}�i-�o�:6^i0����1<�6��_X4��Bm��n�$�iC�n#��T�	�տ�ײ���:�s��O�ڝYk�;�vK+�Q<)L:9�rH���i�]32b�aTJ_MN3����?}ɇ}P�EAڲn_��G	�i���;�"4Hcm�ӈP� �\���"�%��'�fLIŜ�����<�J���<����(�@iqS4�l�G�_�n��"<���w��je�U�Z���X�z0�)M��9��*��7��qv��-8B~B��m�v�\D��bi��u������D����k����:S~pFy
��5�@t%s~}�0�N�@��h#RO�����d�g��uټX/IA��d|赐Nh�b�'��MH������ǵ8: bltψ���u ���4P����f,����Bt���оVG>ͺ�"�^�xK`�4�qU�Ɯ�J�{;f7ΐ �K�R���cU������x/n$!��ɤ�5�Kul�<��d]J7o��Т���(�t���L
���JqO仞��O�=0~y@�MZ6Y=tEA�+κ-�[�v+�������svGu�����ܕ{gͼ�m�����Ya-�#�I�+�H@k�!)�p����:���,f��>�=�0�V�z2�N[�@�+j�Q�$�D���Ueo��d��2
}��;_�<72)��i4lv5_y1�qC���V�+��o�J<��"U�u@��q(��,K�-���seW����?���v-R�� ~g\����;U�0�� �@?d��$|3��c��xb�u�3Lg�����m<7b���^灓�&P��f��m-v���^N���\Q�N]0�pU,�t}��Guݽukbh�`s��e�c:�õ<�N��kJ�~Y��! ?C[���T?[�z���	#������±������B���Ko�$����M|��* |+2�m�#�Oᑫ�}Jd��hD�"���D6�F"a��
W�;m�զL��x�4�J�I�w�^Xȫ*,�AH�P�(1_��~�@�x]D��iU�$�s�yzc��e��j[GfҘ�-�O5tVKs�E��9�{=�@*^It����{U��^m �ʣi�nÚ��Bmv��!���	&4��ܱ�eos��
�D7��ҧ#�+�=�	��T��.M(��袲D�Ǳnjt�<�q�lь�>�5Fm��x����K�w�1�-��ǘKK���9���n�3`n���v,=wB#�[y�c����kX0æ1Lj^��1��3w��f&3}w'na��-n�|b0��3&~�d>zBR�?���!ț����mK�w�L�e|��lT���P	MlQXW ����5\�)�	AY?�O�R�Y�O�^
ʂ�,j�p��i���<������V}py7�e�9-���Q�| [���٨�UsɓҁY�O��m�=H�vp�B)���}}5��	K���>�q�?[���A�bh�m�@4�3;����"�L(��b�e{W����ќ�&��U�o�������Q���_"�F��{��H]����~�X��p�L�Q�qY�.�"D�}}�c���*q����$p&�������T��fH���o��-'z��:Ws�1/Y���i8�lj��޻�q/6jI(`�<ޏ�p��]0�TN�3y
(�Mʓp�tOPC�箖�S���uH�N��4V�>\ˍX�HB,e3���>ʺsp�x��+ł�1)�è��]�ay`�b�Wk"��fd�Z�	]&������;��m8�_��c�J��tg��7O�ώ�0��]���{��/O�ڴ�-��	�[��&��Cmh����]
�OC"ނg���Π�].�`�s�|�A�T����ے�	�:�Kv��w%���0P���B� ��||$й���|���_\i,ѵ.*����s�}��[��*fF_������W���~#�Z��@s$)�Po�}��R�:Yݬtɏ��-�� �{�c�b�n۔u���z�h}��M�O�ϐ�C�>��������_�f,���c�wy�����	��IS��#ߒ�O����>����{���[V1��l���ۡ�í�������J�9j�bU�/��*L�H�0P
V�p󋢯v;{�gyY�;l�~��ZFv(�I1ק!ϫM�o��ӄ�QEk�m�x�	���d�1�6q�yy- u�J���Y#:j��Q�v�Bw��O�q�\�T�w�:��&ֽ���Z���Ю�9�G<��LC1-�'���"o�� 7�ZW3��Ķ��5��ׄ����[vRώ�B�(�� �w��ۜ��C�!A��h��DX3Gǈ3t=��u(�W�Z7�)�t��"��E�w��V� �+��5����^��ȶ�oK{T��@xf�5Y^�����<κ�Ȓ��y�!�#��q�L�
/n48��w�������0.-�6Q9�g_��1�T��T�d���
��ݍ�$>�y���)s<�NZ�	���h�)�˗�%��$e�Viر��oz#�q����nvnޞa$��Q���n��U{ۏ)7��s�VS��@�r{1e0���2-x�<& ��j!�@��\M��]g.�d�Bx�JϺ�Bh#/�	G���K-o�a:��!�wI,~���������K�w�@�?��L���A�E/�p<��{϶^x-�$}'��m��"H�����Z��2>�����Q�)�0�X,�)�B�ErW:�o��5dD��`G��bi�z5/�>d�ϔ�u��|�>vUӳ@x��3�{�_>��:���pFQ�e��=�N�䓒��L5i���ݽ��U�/pgقi��#P�VxW����K�}=Z�,����Cp ��_�(���Me��6BZL�cm�]���� �u/"�3��-���t Z̍�h�4���#ji��v�t�� �~��G p|���<S!��Xl1� @?��ʛ��LWď<W�W�W�,8s���9vN�tQ�@��/n��K�� �c��<4�$����Ve�L�(A�K[�_`u�*��b��u�"Q��x�F={��</ԓ-�5w揓���Q�r:A�D�w�ݤ��.~�H#H�����͈�uj�E5~pnB�s������UKl�(
o��&$�{Ug%�Hҙc�Lw~(_��O|�u䍰R�d���[�++{ؘ��O�� �@���n�*����<Ʈ>2�_���ӱW��o�HfN�;��,p7k�s�`���������:����ѧ��j�/�Q�D���jZ�p�[Es�JA���M�XD�L�5������
�@Jm������y�a�j+�k�q8U�FXj*�-)����wH�r�03�#�H�7L��|��֠&�αn�U����$ԉ���\Qc�^KC��8_�(Q}�ؓ"ަ�C(Ξ�^��"��ٔ�EGςϰ�!vk%[7����=imrQ�>���L�ʹ?!�Pw�j��H8J�0�ؽ��DKP�9�r{}��������U�2��Hx���#�	}nKi�!A0���_Q��@���'�TY�\� uj�Gr�`|���c��e3�Oݡ��;�@��U���T��kN�N�9�����,⚓���M�U
�a�#��K�b<�z�I|���f���/R^D_�?9�
|�MX�A3��C8�k���?B�;V9�a�0��x��0َ%�=>=+��63�3���S��qt>g��+�x��Y%(,�i+�s5K��	Ч�~P���ݻR�ȵ�<�i�gr�fa�i��g+�{�N�δ�N-�I��q�頝>� \]�\;5�u��OY����`8�3g5�;	����oJ��i��8���D�*�z����2Y���n?1���0�y@��P��^��ơ"��~p0z��kݗ���`ѫ<K���Km������f7�� {�M��{��o�����aD
�Z�!;r������8t�	��8z>�*j��������#e�.R[�(��'�.����ь�t�?}ت����}Zb⭕Q�@�K���SzX�3N8�Q:��%GQI��J擉��u*� `��Ќ��~�Q
�#�b��߉5T�-�o�8
7D�n#�{4:��E\�	�X��־;��#:�X�N��(��J��˟�{O�hg/B�De�]�f�=��;E�og�k�H�>' ����IxR0�&*w�ŝ�����#�X��� Q��@Z�tQ �c\;|Rlm9k��~>����]��ն��Ql��%U��vСݱ�e`=�|�e�b�E� �
�i��(�"�$ �������z��jc7l��d�d�����J�?�m��&Vt�����7��oz���[9%��!��c��f f4���-m�E�/�DCڿ{�[��c�k�E;)�WX��Xm���mj��{��3G:��ٹ{�2h �U"�d��	{b�S���N6��	h��+b�*�PP�W]ԕf�-��)��eX�e��o�T觟��O��.�hx�;����w�f��h�>�h��܏Y0D� �Xk-���yY�/<R�GKw!����������\����Tn�I���<S�-�	�7�sU6ֆ'�+��*���4"xE��`��J$k����~�C
$
���K[)��bD5��UV������*��faD��
���\�6?�������=l���`z�<S��y�u�h�����>����D}���d�r"F�;�O&�0xRx1�au^���ʹ�`�j;e���%�z�K<H�D�2���{wco{��Bs�J��5�Bx�:����ym�:σIB/'7K�C�P���U�
i�!��<S�1a��\�<�Q��Fe���b͖p�bK��	���,�*1�7/�zUOz�5Z\�	�%\��J��vK��t���臛��Ԫ5]$�h���YT���?e�J`���]��q$,VeZ��a8������32q�=�,g�gd��fwKN��6΃���Mh7�$g�aY�\@��Ut���GG~F�?{��/m�Q�O��}�0G*̃~|U�Cn�w�IW$���1����F�!+6�XF"4F��
X�g��8qc�����n�u�=�$�"�;Z>B�kyW*tYs�)������!d Q�:�i�4�V��J�'��H�Q`�Jp2l��]�Z�Z*)f�[��M���nyK�o�3I*�-Va� ��c�B9�ݴ��q6�X���Й�	.�:$F$S�����e+��T�XF:ا���-�Bs*��M�U�����o����q��S� �� � *I=n��V8�R#]dl�rs�m	y�-�6�>*qN阝H�m��P�m��8{�������u�[�1s���*��Z�fv���������V���7��}����OBA���Qs>}g��>�	Jv�x�y@ǻ#��_���"�-̱� �a5��o�
RJUrf�2?_�����
Z�ݛ� {��?L^#0��e�_6%H��Eb]L����0q�E�L]��T�,q/��Y�ԓ��(��钫�bQf�;}A�����kjpP,쵏���`!m׊��/���
���2Q������u���Ã��yKE����P>A�THH�&����Al��*�ͺ���x��+K
,���=�nu�=���f�\���^c��V�Zӛ�����{�MaL�!�~����N�DGH�����B�]I�F9������Xh��՜pL:z��F�{.'޶]ԛ�Yh���9f�i~ �O�G,>=L������,�R����j��!�2���nf��^�ę59��٧�,�(B�;����
�!n��'+�Ɉ���sR�''�����3r��{e��?����մ()])=��Ƞh���#��Ϧ�ru�{Y	6�u�T��EfB�|�ن�֒�p!jZ4k�m����	K�� �~v��J/�����e�_���M�mb�b&��:�&C�<O�G�� AZ�G�݂
ds]���L�� ?B�mn����=v�4a��C��&�q
Dd ��?	{H(~�SY�?�t[|��xw{e�2�'2�7ĝ�0Cx�E�7��W��7�����wäA�ǡEn�Gq�Sp7L�Z��q;!����?՝ϪǾ��w�TW�(/��ڳ�s�J�C��(�ٶ����d؛�Ҟp%us^��G�2?�h]ƨT1���44�z�#\WN1c���t!l#<��7��mX���?uȚ�+hMl���3�v��$y# HS֢��d�� sm9�11"��Egn���}��z��]�=���g��`DDݤ�X�A+��e0}�m/$��F�tk�X�pXU-�=�p���%��JG�������K�NGo:ҁ����0��)��ߠ�hGM�#^�D�nThbJ�;ER�S��h�[N�����4t��1��R��7��@P4�U�y'F�*?�D�A�����S̧ ��ar�v�П+��NdzV��$2��ť|I F��\H�/LYŐ���}6���9��öJ�J��BA��c�t�F�C�(�����x��$ss����2\tvM�o�9��΋��hEX�&V����~	ꆹ�QQ�W�\ 뽘����Bh�@O�����~3�\
�d ;s�ːf��{��C����!*1N�'o�Ne��T��QTYn�TY�mh��Ք[�C�_�o�����z�ޔ=�$�������Ktl�7#�����Oz���ךf0��\4��F�]�Sk1���X�&�(��Z���S��^����{lF2��!+B�RZW7�O
去ʊ��;��zH�(�8���"�&��Q[��>�8����[�{!]�e.���ٴ#iB�y�[�8Y�C���o�nb1+�H�YC���5B87�T�+صi��5�1�%�28�.�6�Q�拗U�i�,e��Z��}�$.���3���q�i�~8xF?��Res�-N�Y����"*F>��{���[%g����Kr�B��W]�����U�?����@��5�aV3��V�̗�'��p�Wb���|p��sP,�Y�6�v�WB��Xkf�Ϫ��s�T��N��r�&�vA�l�l�t�|��5lW�Ȑ���[�Q�jK�77�|��6H������3������4m��d�W���xK1	!6F����c@�1�\�9�[_�NE�E���p��Ɓ��yOt�������өM6K	Ώc"S��
��]:NN�1�jK'gF;�X�ۡ
�ڔ2c�㔌��Sn� �­
g���=;�`0�u�c=iq��P�v�K�7��P]V���}S�R����.��
���d,
>�9��L�R�/#�}sN����z����2D��;.�Dr�gA\tS�f)=�r���cFApͺ�z��Ǿ'ΐ�l�n��B9	؛lɇi�;���s���ײ��p}4#�Vm��ZJx�JuH��3�#E?�W�J����ig�S��C3�����^��HT45�G|�	�8�߬J�Я���,e:�1�}oȧ�H�+�;|�d����n�$�~�|4`��n��&p��/b����B8�bq�s!>����ab'���0�0U���"������h����l:z0�1���������y'�88�S-�i����0�6-T����\?��94���+�W��O�V�:a�m����l���F�b;��W��Ɏe�n��{��Ϝ�(�u����Et�1� ���VA8�l�U�L�$-Μ�|��89���{����q��=j֍��W"9j�U���3~��W(_�[a�.��E�r"�@r\2
mL`�ׅMB������0���!���(�/j@.!�1�ĳ�̈́zfA��h(Vt�3ᣙќ���&��9wwI�3�h(B_����7m�����P[���u�/qs&"qAO�5��{ /��oϼI�;s�f;#`���[���İCZ��Y��QjA����S�´3�XDKS��ټ��赛a#Y�>�0�9��!�{ز
�؃���Zg��.Z&s"i��]���0z��`Qb y�L:�3���pV���3��Q\/Y	<�>��u}�%_ �a42����L"S�+�{#�"1�+����,XX'���F�F��V�#򹮁Wa�����>[H�j���+_w�]Ҟ���m��c������)ǁ�wp�)�@ ]���/e���E�B]����%�}#��4���eQO�A<D�m�4�(�^������F��1�D�vX�؎Vתs_��#0�[6��];�_p��O�i���>�T�:��a�C��$�� _Gf�ev'd��RR���LdAR1从LI$�ץpØ���6d�b��(��F��)9�ͩz�J��oI��	!�� ��2<��@9�Z�vS¦�\�E���^��}g{@�X��;�t@W*u��*tk��*\�]^ Mk/@NSz�e;'�%�ƪ�w��O{D.�T[	W>���V���G0|���ظ��GDR���d������%���D��ؠ�(�ޖ��U��z+�195/&#P�U�Xu�?1/��%����Weaf4�g�/��Z�<?�r%Ơ{b���$ޙ���s���h�_.M����H�*Q���J�$���a�܃y>��$�Z��/�皍C';u�Tѣ\ ���0�0C'O����[�ɮ򠸆;�O�;�F2��*��s���.��5Wc�m��a�O�s��6Q��Vja���0N^�+�AW��k���"��g(ۃRa�*���U#ڄ�MH~Z�ѽp{�,2[2bS�a�Ő����+���0��~Ӧ*�)i��k�^a���P� $�#hN�ZA�[Q7P`�(���*�zm��	(YH���R�Y���)T�	�v��E��fd}��޺�����u�̖�z�sp�'�6�RVtS(���0L[�������ga�"�$�%��DX�ߙ�l�-,k�յp)�C�=G! /���6f�|��:�Վ�K`4O�B�%�Z2}��b-ͳ�s��0�\JS}�;
X���V�H�{Aj�B���GG��"�����YN����}�i��]�Y�3������ɣ3�x@�Uo/,���$]ޣ9%5.�����X�_Ѫm�ܧfN;H�7#�vKl�'^��R���0ꖏف𨝼��2�F�N��q��qEB�n���U;-u�%�����䑊*����k�c_��	�[\�B����a|�s����:�,�.M����ϊ�z@�.:���E�>�'�ߢ&���4�;L�;��7��jZ�n�� ;�M�C5JQr��Ũ�3G��p�|k�Q�+��.���ip�o6�'%��a��y<�R~�E칁85�1�X_3���Y��������P����z��[)P�
m8���s|���Vw�A���UH�_�:����M1���.�
�A�S��X��I��rq[�iA�'r��v�>Ez�ZK���B�ikS~�}H�R����{�#\Yc���z����_����9�M%d�	$L�����=Ǫ^*O�z�a	�ޟ!����K����9�(o�K��q/�W�#� X�T�O��T�<_;�t�ߩ�;!UG�ў��0�efY��Ȑ���PCM!�:�y�C�d���+Z7�w�i:J�Yz#�g*��q�?ŋrm���MmZd&_�N��S��_;�ج�8������{��q%�����?ӑڄ��ąk��?��9��W�M���O}?���!���5���g�Y�Jx�k�L�X�`��[|�J�Kx8i�Zh��>ν�q1]6k���o�/E)F�>:c�t1�t��Qe�VwV��Y�޶̴G1�ZTR�Q�U%��̈́�	y���}Qe�!=�3�|e[�wM ����J�n���M�[��X�fz8�t�k�G!Z��$7M)0-jk!�^�rz��ɪ脥��1�[
G! ���|�2��Kq�6���ӕ������U㓬ȑ�b4u��E�<��I{/Ƥ�H�?	��*������[�|r-�>�n'�
���7�'���o�F�bJ��5Q���^���R۩j.|�V]"��5�B0�+�
��s�C���c�x�`�Zk�;��EWB�=�����VR����~|S9��SktKo��%z<�8��F����W��n�?�,��m��e.q�]TK��.X�u�d�����
�y6��(*:X˲���$$�uƽ�
��M�.���y?M� �)�B�¯�\kaf�?�T#�(�E#�_�"��'�UJ7a݌�ǬF,otP��l�蚳��|�3H�K!�Ns;�-";5���8�1X���&��6N�th�|(:#��?Xoc�[��/�B)4۾>���P��Do�Y��A �E9��\YVa�dI���3E>x�g��3�'S������aՎ���H����1�(��*:�[~����?�#���
R�������d��z"��4�y�������ej�J��a�O��O����{�XT�R6�l�������{؜Mc8�9FZ��1������� �Oe��]i�fB���]�E8���>��f^F��Kk���>��X��*��)��^��^�h%���L�*���,�>��[������k@��`�
��V�z�6�>�ɭ��ݬ�SWY@����d�*�s�Y������ӕc5C� ��rxj��9�^����D�x[i,	��ޙ5�<7��+��`�܄����N09����ua�]�A(������9��N��І��њL\H=��ܘ��H�j OA�L�
���]�u�����w!����V���AѽH��=�ݢx���;	��󊽫mVH�l�ზ�m,=v`�6���`7�|)N0 |%ޏ�8���H	�>+q�"�:�|��T`�4���S3-U��nB�{�_�~۝��/�� �����^��B�s$�ک��ـ�9��P T@�����6�]=������<����N���7J}Rm�������V�ְ�ִy�x����(�ϭ���D�s���Mi�2�`��D 9�O�O���)��Q��4�3#h��U�.�<�[/1��a\�� `�pR3��2�1�_SkB�ݎ�ITKQ��0�3��G�͌��F��n�G硑~��ݜP�6���0�D�!��.(��m
�Ka)�K9e[~R���?�x�����F�M�;������@$�c���7piB����J$�)��~�yX1�==D��*(����9H�����l����L\�~�?������ଧq��I}!R(�˄�#�uZ�ꨞ�~k����.a����V�́]~���0�r���ZTY�������M:��gi��J:���Ω���\_����Z�4���6!=��6V���=�W����L%��"n��d�� �V��(|rϙ�o%T~� �Ni:'8�� .xӄ�+�)%�M��j1?u�� 6x��rƅ*(�V��6�	�R�b��������@����d���/�#�3�[i�/:���tM=�S��ԝAw���0������os#�Ȱ:J���D"R"�ڪ�7���~���7��sO�p��O@��a��|Q�e�WI�u����+��Yڤ&n���0B+x3����Na5��m�8+)�����5F�u��}6!����#��"#��n�6x�zJD8��x�CP9ZW�������bN����[�.*�Y<��"b��x��H��2ڭ+p���6���~V�B��h�$$�a�i�>��JY��>cқ�*<=A��E�]@�I5�����Y]G��ѭLö�>%a0��Ƭ�֕����������P4u�(\�#�a:.�jI��"J}w��$�'�ތ�������������0c��1��H�g5Vo�����%�9>-?�W~�W��VFT����
]x`_#/C�(�XT�0]���N_7L^�̝r���`��	rd<�	�W����~�K��?m^��y�?(&���ᆎ�̴r��Ѡ����ԻQ�d\�	�Hd���㑠�M^\�);�ݿ3Z�ȅ��z�fʶb�=l鎜���v�����ʃ_X���%�G�6��e�b"^��Ɔ4�}�(���,>���8:�?ʮ�A�*���8m}Ҝ��骜�k({���qG���tk�f*o���p��Ԉ�ڈ�߽r�����v��~M�R�ao]
�i�U䶻�p�pO'<W���_�i����ϓ�AF�^d��0�����l�/h_��b!�ef&�t�Iu_��qrK�9fԉAѠ�S���%���b'�f�5pD����y���0%�l�p�n��� �������p�Ӂ;����T�Vw���
H�p����P�h�m#A<頬�~Ѝ߱z��Kcq�;�� �Q�0��^��ǈ+��h%����c�Re*�O ��y@�b�qAdZY�܋ק}��X���VY�D�y�kN�%R���f|��R/f��{(
��K!s/��A�ݟ�,�f�u�9���������V ��2��D�$��nU���z=Ŭ����`ro���<pRQ��&���:��wh��E�:�'x�uKV_y.���B!�d�	Q����\Ұt�i˯Z:���.�A6�^����f7\M����83�p�"�҄���k1�wx�X��5Q��G�<gO=��Y{O��o��MDk�p?����w�n��_05 6��.�g��Ԭ��̘QV��v��a:џ�d*�S�q3����gSK�m��13�癶&��
k����@	Ʃ�C*���6��˔�>�`g��;T���]ȑP���D0DS��ϭ6�d�ǜ��������ZX���>:1�N�X�yi��S��)}�����n,�	]�ҩF��GgT?���>�t��<l!����y�@�zY:�¨�Y��X
�g+ga�	����:JY�ӷN��*�]Om?W��t�/�as�Ҙ��o�S �{��r�}y,q�v�>6 
�N�$P�������Od����[a�f��p$^��S�cTz�0��#]k��i|»�N���8V�Xsa<U�V)	���X�!���?1}t��wx[�թ L�F�-KJ!-���I�͛���8d��'yzE]�{�?���֋S�|7����Z�w�m}���x�/��Dށ^�=�u+�dE���>��;���rܻRz��[ȫ���8�CFϼ�=�uI��t��)��(�e���Z�ղ��ôa�>�M�:�=�&�cw EE����d#�7@z��.���v��k�I���.�E���k:�!>�u2DI�`�7��a���
��o�4e)hh�dބ�y��N���=ڀWi�ʇt|L>\"h�։8;e�5�˓k)�6D<� �b�=�si�Ju��qE*&o ��m�B�ߏ�3�!�+$e���O�,4��W]x+�T�BY0�� �]Sy�0g���Xć Qk&��e�� u��'���y� �Z��^�u�+#�d�s1*R�$OĖ�1����89b=oCAjJ8����[�DTϷ��s\��,T���I7u���ĵ��=�˭�N�'g㝹:�o;�������NPdrs��P��͕mϡ�Z�P���h�L�H��+���R@1M��q{/�(��)�����۪p���˟Dl@ȳ��ER�.��L�t4 �M�%~����/S��K��I�W����	�d-	��w,��-�fw�6���:�֓���Ewv�4����.>f�"��#}�f���Š{i�:q�J���&ʎZ젺��X_C�}�9hr����&[��0�+�������j&b����8�r��UWnBA��e�ҋ�'Y�\�������Q3k�m�3��)j��0���<�z����F�b��%'l���ٹ���Q�� z�e�leZ(��aL�Es�⠒G˳/<��-��C1�Ѵ~EV0f��,���pP���i�������so���G$�s~m�M�ذ�U=�׃�R�jt��f�~���J�Z#�󽠒k�D�x��nz*��~lo,�c9�m5홞�Z���@OsB=��@�����9�P��G�Eb!�4���$��D' 0�j'2)(k#8��뿝�w�8pk!��r��+{h� s�DT���F"��������*����d����[�0�X^Jr��f 6ȸ��x��:-�����3cQ��p	��G�O�02��L���u�U>u�:�RP-·�[���/���>&�"�v����S�	ߘd�0�.*pӣ�
D+Sof	m388GHW8�R��N���}�ʠ j�ϣa�E�H���Jb���CT&.-Y�x���|�@��Q��6����)*�B:>R�{fb�����_�=u����Ѧ]%o:&�̡�Tb�' �̙곏zoC�㫥�57:On5��"��r���%%������r�Z�Z�s?8���U��﴾eg'� 72��BȽ�)��]�+�H�a�H��[����m+8�E��XKР�m�4l�-̊y�Xk�2"�ܾ~lOB7��a��b�P�\P|�7l%̴�Ȕݡw�ʇ���ο�����6��j���ԟ���`�� G�\�D3���CTYfA9���i�V�A� ^3W��L?I]�1��^D^�2�q!��qb�v�;%�p�t�L*��hi�����G�"a��nkr5Bwg���؂(�'���&�ܒ�L_6r8�nVt������u�m�񉾛�qP�9��Gg���§��|,�~#2��6� ��
ãv��J���/ƙ�����˖�jhBD�m�d|��4��>�|'b��O����� B��BesG�~�X8y�'�g����j\��	��P}4���s��'ؐgm_���� =&��ax���k���~e�ё�>�=U'	�FF�݊P�L��e��XT>�nǲ��T���T�(� R��	��<�`@(NI��f����{�"���v�~�`�ٗ��0 O8��� ��W�U� ���kk�����GM�e�<N�@�H�A79�"H�)J��Hv?��y�;U.�奍���ծ��:MӃ��VQ�|Y�Li��Sӝ�EQ����S�9����G|2#'�.�0��,�J�P�=A�½8�T��p�	���n��{��`�U���VF)��*�7�,^��r^'9fx_�|�$��\�N�_���XD�ta~ ̓� js{���*hW�oթBt$Ν���aw@u������H���b��яF� e�Ua��S���l$�L���� �^���+ѫ��h vB'Ŝ�#�"7�ʰ^z�*��4,y�>�[�8S��T��쳺ᱤ�˒��4
�8��pZ6J�d�>���F.A�!������mUo�}U�w~������r�n�Hܵ7��K�pXN�P�z����8�L6�t��.ɘ���0�#h�I(s����T�F@U�qQ�va��h�Y��t=��ds� �c8�K�+:��5���>�Ç����t*3�h��D`7ۊ�&�*��gf��]w;��"p,�D�\�~[K�2 z�C�x<!�B9�*b�����W ����yy��^��YS[/K\�����j�1B[{��p��Z�]$3u�|3��dHbÃH!�z������Qr�׼���K�������]�;]Kb������_���NO_����W�a��xZ�oʹ�J�VjTY���c!	��@��y�qԞS!\=ŢS�}��(0�B�Z"�%��7	G�&��F��)��!����<qRE�N����!H��K�����C7Ol6�M۾2M@����j�=>?g���@l�C�Q&|ڥE����F(:X�s�T~�$�1 ��L1�?�ʗ� H_g�t��ɁB� m�@$��HȊ4Kҍ5b�l�G���ώӞ6H����ekr'���O��}��:X�/#�%�%1��WEz�?:�I��c���� V���RN	ӝ6�'3�x5��]L.�5��[�c�$u�
������1�#����+�=T��k�@����׽�.9���i�j���5f����Kˁ�oʭ�-fPt^�!L��HBQ�̃��k[U�s6�wƨy�v��S��|���|�.�>X�.Էu�TG��-�f&��Pu�r���:>S����L�}����P�W�7�8�U-��(�؉
�)m�U�ݢ�\8a.��T� ��	�IX&�����V`��	���`�k�ÿ*;�g|k���oc�M���J�3�������n�:~������I��o�KE}�LRyU�p4���1���D�ɇM�Y;8\�����U�}���5�q�˓HX��q1�~�d�h���w��ж���0�ֻ�k��}�3���Fo�1G;�G1KZ.��T���\���7��;k�Ξ��%�������(�L�)�J��#mߧ���+=a7�z8ϩy��D5;�<;��Lڳ3�6��I�����wq�2p��W�d0D��~?�4�w$�݌�KmhJ1�B�<�A�5��_qWӚyN��9�gQ��s��1�e��6�Բ�������o?��D����fXGe��di��}"&��Q���טIR��C`0E9?�%E��� 	��d��z��S���P�n��W�]���@,��;��gs��[�NF���Mɹ�A���}��N{������أ�H�rܑ�8gZ�T�HɃ����	H	��*������,��� ��y4��$ AG�1��c�����@�31��R0��)�Y�9���d�6�����R�O�����Pԏ�RnM�����04�[�Y
co�u��8Ac��#f�&C��gZ����������	QW}����ˤDÀ?X�NS{��r�"�d`�$x�י<�O�.����[��5T�(�A~<F�~��u��X���Q����>~��u�![(����$/� ��Eo^�M���ϳ��=v\��Z��a�����^�2֤|a*o������r��Js]uDⴎ�Yп��?΂<�G�[մ���?N)���l-ٞ�j�>��Ʊ�Sԁ�r5����D=ҵ[� a�R���p����h���������Ŭ�1�7Y Ԟ��a�Ϳ��ڌ� �_p��s��}�+z�D���XF�S8@��9Y�h�RQ���ì��~a> �YKj�eFxJ��s�Q�'vi�Mn���ϣ��ax�;�D'�ʰ|R+��I�$>:���Kb��F5�-��bK���.���H�A��[��_��VS�a����Z'�~qf���*��%HH���b�2��:l�kǬO��&������̆x0��Gc�Ne����s�e�p��;��cGiw%�$g5�A�V�c��2��_�,\y������bބ�R�y����T�-�z�Q���Y)"�t8m$g1|�"e�(:�!�Z�������]�$��z�o}���ePb��Ἕ�ߟ�Ǟ>��x��ss����?�o|�Ra��b"�14,�4���iA�(�?p���L U$�.������粑���jAZ�m>����"��C�1�H`_�,��9B`L��#�NU�p�
�Q��.����A�#�D5�)��O˔!�8�;�l� �N�{#��v
���#\�NA��s��ǨA�
�s���A�:��"g�*�����D���l��K
#lg+ !�9���� ps�+�=�n�m��GO�~�l�|��j��i�B�	F��.#�9ޫ�NFy�cY��%i�k nljT�^W�1'���F���)�	r��Ҽ���F 0�~�:!�� DC���v9�_ЋF���/����HRb���K�v�*T���:�ݸ��V�����zjs�Ԧ�ɘ���vi��E���}���S�����BG�-5�Xes�~(+���s�擿�bMc7���Ԟnfg5,��k��6;�m�: ��*D1rJ����DI�07�m�M�G���!�EA��;":j�Z�8����Ӣ�J�c1�j����W��~�M���O��Ü;�����h~�����&zK�t�s���ay�D�	��0���"�=�ٰ�yƇ�����adt�\8����k�w�oz;�i�HG�������σ=rj:auc|�S�� ��0b���]O�L��[�T��=��2�f$@�u�����1�$O!(������&�(7I*��5;�/��s��NB4��iS�Śɖt��^:o�,8<U�3��DݫPѫ-�-C�	o]a��BRDV��5AsSq@'�� ��w0�\��m��t.�"����tf3�op�>*�E���� }d�{�tP3D�Ϧ���Z=�)H�YV5��c��Ҭ\�[���W٦.���r<�(���/2Ь"FXd$�ʴ;Y.//xy��!���<G6ڈ�Y�9�x�Ȏܿ���?q�Z���U�l��)GZc=�;�e�m���>���&�YnE�8�:�'i��;��=	\;�#Pi�'�oqtr���s�,�~���k4V�5ei8�̬xq�3 �xTH�G>�������3^6�"��ʃdR4M��C��������N�%j�����2ߕ��Q�"'\�^q�#��F��z,�k���{��d��>��F�6>����a|��vxf�RiT�8O7p���e~ji�hz����_g�$�y���|�<��W]Ҥ���_,��XB6��e�n�]�`�n�F~�M$�����ʞ����h�qiu��M��d�:-���ߖѺп#�'�s�OeOZ�,�POw�5�Wli0���z�U��*j߷�;z��� �B2�3�(�$krp��S<p>P
Ic���H�"�-,b�a���9R|N�Q�3�����:74�}��o��+�5ܭ*���yެ�G-4j�.���2fk��jg	q*�Й0�Ͽ�Uv[�G
�;E�3����˅�`D�e~� ������q���M�I�6>�V?�U���e�4Wɶ̈́�\O�w���RF� �yQ4���,ɦgRZg�j3�Ix2%1�D���.Q���5���Pv���0� rH��E�<��3�+��4d�o�b;K������5ڸ����p��%����5�L�����̭�e2��	]���3��ծ�����ϯ7���,E�EQ�}cVΌ��r��,��4���`Ħ'Z�������Bcf���[�fU�`=���T2�>y�|�e��?��ؙ�ޗ�[�����LW�%L����}x}�l 0��<S\Q�Zͯ��bJ�ţ�?�R�G�Ӳ3�j��@�:�\�c(���$�l
CW�x6�fxuv���;�/�o�zFٹP)������>.�=���r�v��4��~�,���jv�Ѱi�:��&���F���t�w�H���_#�d;a{��=�K0G�k��i�qM�ǉ%2�p�wk&X��R� sE��U�C��ɢ��X]�)����k��4���=�
m�\�:�_��Gt�k+�q�B�׻��Fw&�B�@S��z���#���Ef/���
�y��ZBŋ�;�b�E=�>���vv����S,vJ[6�:�6.�kEV�E�b�+�6 �#�ĳ�����3��`�F6�)sx���;L�m���;?O-"�j�ɷ���*����-�?�D�1�(�I�G^��خ�k�J�1���YIQ�*\W�.?��~gJ���7pob��P�1���"��/����_�.���̤^�$�U�s�w����4��pyXt�@�O����_���={����4�[v@M���3F�����u6��?���i~��8p�;��o�$k[^aa���R�f�^�>����*hx0��hNJ6��R���5� �uA��#�˨Ǟ�Ddީ��ha���w`����_'vӌi1GT��MA;�w��)��E��BF��?��3��-hz�|�UA�"H됴 L���nf�3�mr�3�Hl����6�4�{A � ���A�>�IaKc��� X��7�?�	Cn�ǃ��Q`Y)��S���B}r�>�2u@�]�?���j茮�����$M�n��N��˨4��%��J]S��oU��*(�����|�a��l��N>�ͱ�)i���#4ٯg�(j%��F!W��Oƽ*4>U<:{�R(���Z�?���B2���ǘ7e&�X�v�X�ǃ��[𭈭��gb����ܸoJרm5/Fȋ����vz�2�Ѵ
���|��|f֊�B��ʢ9� o�3���I�� *O9tjc�O1q;ۻ�y�߅�:X��$6bP_xQ���e�6m��B��В��;�e�7L�]D�c�Wr��/2m잤Y8�u��íe�ku�70������0j_��r/�Cs2����F�-���Q�!\#���� 	�����P�S�2�h������I2s'Q� Y����]>}���{g����7�QJ����vx���=N}�;m���Z~��z�-p�s��5�oLA�=i8bW��A�Fi�	��4�H�T9�a~6}�@�_!x���bc�I l��ƿ�*j;������l�I����0M�%���ɥ� ca�ؽ���8K<�J�=��������9ۀ(�9�`K�^)Cy;i�=��d
�$a'�D�]N�~r��wZU�qB����LW�dee�^��V��Dr�3�/@K	�o�3�B�v[�9�՞pp#���[���u��e��۹\�-6�A�|�0�� ��<����A�:��?
�7g9	�l��Mos�pr�UX~v�V�t{OT�;c�u��{�"W�k';e7��t �uOxyxm�!��O�l�J��$\�L��!��IZf��$����
d�>�?x�"���eWa��/Xb$v>���[���~��X�����|"u�ʿ��[���jd9���5��c7w^b{f:h'oHn��>V�"g�|�J����Nƽ~�i�$����k#ѷ�p��P�������<�*t�c�Rn����"���P7ZKۂ���;t��`8��߬W��E�_� �5�5�&x���/3I���7�"��ǿJ�Жs|�sC�E�|aE�g$��[�g�On���C����\�d��#�5��G�k��>�מƛJ�ՄA,g����E�_#iܴe��g�+j��1�#�a���׾�f��S����U&�?���g9�]�Ꚇ[�9%�����
� ChE?���Z
�پ�����a���0��UI�]����8b*КC�Tl�'��I)�i�_��w��P8�����xh�Hz�r!;�����⦪�m�
m��KB�r+�ĹÓ��@����z��wt�?oF���,�ZL��ШJt��i0�<�69	ϐ�fV#�y��}-���pe����_C~Iݺ��(M1#+^YcP�k~e������/�+�P�ch�Jm�#����z�=�	S�[��t�� ���B�������37$"�(�
G��D�mwMr6�l��u+�	�?��U
�Q���'�&�X_�A���u�}誁pp:�������������Y�`��Q�x�Td0��r�I�A�;c�7��5�
4dDw���BN���(_l����R�m�{R�>F�Ņ��h�}�w$C��ҚBX�W3֞(es�.���B#S h~/�8����!��R�y���ʬ�[VYT^��sR �l�f�{t܄xoa�=GA,��>9��w���DX���&�1^�e�%���h_���z��ک�.�n1���w���c$zJO��A%�Si�d7akͮ��=K��.�u�/? &�i	��,y�y*��?y�W$ϵBb���`8))�];\x��{��e�%���5͘�#��l��X�@���z��1������u�y�b���M��|%ѕ��>��+�J�s�{gA�^Fdm*n=u8����O�z��C�7� Ȳ$#�?�֜YH>�5��:�z1Bgjܮ�`[�٣�b�d�����_$��G�����K�f_�n�m1�����iV���&QC����,��-�!��ߊ$r����z��z�/�y ���H6����j�ۥ�� ����1>�d��z��Ie-޷�zZ��i����,˨qnQ?��1�R��(�1g0Y8>�h�Tr�P@�@
�+(Ϫx����ڥb�\Ǔ����gŀ�.�J_و4���1���"�2�p��#�ӏ�e8�;�l�6F��#8I��	��H�}o�&���в�P<[���8���=?m���wԝ�܇/n�'��nF�״��+���e���)�Wj`����Dz����ذ.�l�0 I��oD��r��*��R7�FV�l�|����z�T;&��+m��SD��ٗ��8�RŇIs!�l'
�b� ����=wv�;�ʸ�hoϛRφq��b(|�06���Ici?���!�gBC۾:�����d�� ��&[��Qo�I'����#�=�~t�-|J���z&D�m��#��%��ŹY����8�x���	�ۖ՟4����xj�7D-a�����oy������m��l������|�&�3�AK���s�Nq�N3�ZJ��R�zo�o԰0�	�o�����
B��S�	��ȓ��@+�a���)\��c6[�Ǽ�C�+�`d,Z�=+��s2����Ƭ2��*��r�?�Rw3TB�x����+��苲+й�4Mm�$����9?����r%�� �wreC�A�n���!�L����;�#�!*�u,Ǉ��Ib���t�q�/�O	��;����oSaL�P�iWNz�Z�(VK��H<M��y�d������s(��0����#Ɉ��҂j@N�sTB����@"��0+������������j���X�@����BO	�R/M�Qͅ�Ma8���������+�����W��
�1�c�T)=@[P���g��^(�@�:�Yנ���̄*տA������ҽT�"ce3���Yn��I(�'��_��Q���ca���Wf�5��J<��+��+ �Bb��H���,ܷ�� ��H�,@@s�J�N�|c�g����S��י�=�%�(Y�&,Q��Xj���H�J��;ECʧ"m�V	�}i{�}}P�t �AVF�b��)1y�^��rZDx�NFs�KA�dno;�.�ײ��oI*� ~9�$�8�'���U6���(�f�ٵ������y#@�Y9��1�E�+0����������W����O�5]QՇ%�X�B��.�֖��3's�����B� [��ja޵"����Y�����?B���,��5��(kV�]�S���tb���x��or	^+h㜈�*���}�:���!�ȡ\m��!���1��s��r�G2c�˺�h�L�"^h��>��F�������O9税]�3�~��ҋ��6�L"�w�f��G��;*s��O�
�׉5����Ǟ>���	0\/q'�m_��IΔ~�=s��2n�36#l�,y��M�Hd'��� �bᇼg{4����b}5�H/��ځzYCr�S��[�����~�E�W*�^p7��v.�e,צ �� �A�ጣ�)�!�R[���y��Qc~�����].�*;�r��.������|�5������d �^����qJڰc�t����HW,�nچد�~\�Y��X&����.��Iyp�9w�V�n:c(=�D�c�awV�5�l��;mg�D���E�\H���&gZ�g��2�>3$�z�hV�G�=�3=-;�,e�Jz*m@@��"�0G9�.^Q^_砗��g�8�J
�i$�M?���'V&��U4��뜟�DW<��y� kY�etX����������Jqn��P#-��yX����}�ҽ�$�{���(0}�
�z5r��U�>�Au�=mi�<G�o�6�h�i7��Q> iZ��' ������N���[�6?��ئ�e�!S��L+R�.��I��0���{��9�ב�:J�7wZks�v��>�ۅ=��Y!8�����WT�ϞF�_�(؈aSi��[~G�s��>%�;��&ܲ��W�dz�Þ�urg�$5�Kwuk?4�pY�7�'��U�z�k5���%���3r"d��IN�����7Ne�܁�S��1���oF�\Y��o���CYh��c��F=�h$.�כ�9�朵1yn ܓ�d�ix��!�:�*�۶c�<��Lt�N� ؍T��/s���wS���C}�++�!�S����&s�D�)��@��n��ޙ�8���:��G���Ќ,��Qo��K]|�2���:�6Mo���z>_�JG5i�Qa�Vx�&�2�u��N@٢Rgu��\�O7h�r}X�H�r�U uX�6%=��_�xLc�B�&�2#O�a�@��l��.7y�G[���,���O�����-h���q0�˙�(1�\�nfar�f�^�He����"�9�5���|q�Ҹ�q��X0k�P���F�X�#����f9�2Gp�zH�jc�Uљ2�,��צ����n���J������I��6��yQ�i�R��x� l���
5�7�Ƶ����|C���_�b��;R��>U��ca���'���mLB&���]���V
�3	5 s]C���X
}��P�T��=� 轺���Vt�z�|�kY5H&q6q�W��"m������&�x}�h`�;�2S�����q?L�_�GS�9��-\wUa��s`T�\�ѯg���������9�Z���5<��J��i�.���-�R�G1)��ԃq�[���)32S�NN��zg(�r��jL��UdH>� M��c[Nɀ񘾸 S�&�\	������톭VL
*%���!���_�b�_0�\�J�V{#�����v�m��5N��:�ȵ�~���#�5�$�iB-�����^a�m��8�A�m����fՄ<�fo& ��l� �X�Z�2z��3�z�$�i��ѳ����
\���p��l@�.�
�� ,�R�*/C:��U� z\E,��z�k�"��
F�?����Mi)�����Qq����̊� �hi���\���LLm��
_�?�ȳ�%�*�텖&�³�ȍ0,"�e�Щ��ŵs��2��C�����:
Ѳ��Ե��{}ɩ����rPE�*��!n��G���
��BSRA����Q��������5�w*`]���ϩC�A1[lÏ����r.�1��nХߤTy��gmF-q)_���ϡ�:�NF������j�$�b-�@$�S�'��9�u1jy�s�LԘ��#�ZmG��dR=RKr�m�bG��>=U]v�j��#��y��`�Ӥ�?��f�r�?�j��@ok�D��lz�W�j~6�A|:D�D5�I���?R>���S�*?�@�Dk�OE酋4d�Y�R>a,�w��|=B�`��I^�M�~���*����¸d��Y"�Ug�B�÷������:-��t��S'�Ne�*�;��\5s�����[a����>��o��ސ�de5z�P$0bo?��m�+]6¿e������>͑��M	��/�S�T�vۅ-�M�{���~�
i.�h��$Ł/D�+��1�{>0n/xIǄ�ޑ�$�}��1O�ɍxK�I�3�r��֤��7����7����O���4j������p��x��

8��y�G��E;�E�¬��L#��=��zhF/�1�-�!��)]����&�NP�H�}nB��q:K�m�[;�@1|�%A�]�)���:$3z�%�7`F��+����ri�]��܍��XcA� �t�]B�k�6R͍�f�1��0S ��q^Љ��]�L���.*��O���z�zwl��g[Ӫ�����9Y����J0X��Mœ���`�D.�&-�����d!�iQ7�Ѻ���,��^'.�W0%���?���$���6í|'̀�ũ21��m�&���"y���|�.���s�J眚�$�UAMl^o��!X4��a�Wv����m�5�ۿڬ�Ț�'��Hd���p������y@���Ǹ�R�OP�_�~�m���N��#�/��,���Y|[�Bz���Ǜ������[�Rq�=	��-eEx_,8_���Ch'��v��J�-������a������"�V2��c*�YT�@�1���y�<����17=E���2x5:7�Z�e����[1~	ɸu��<{��GN��-�Du�-���r�f�!���4��k���X�US���Lq_��
�,XsYxm.�"$X9I���zDp�9��ҳft��#��͢v~���^���>��e������Y���M\��/sK@�b�ql��_�[(��۬�&?\��S�W?���¶������0>��rF��-�
��W�����@�7��|9���PO��ڥ���7� Z9疳<J�3Pn�v��!E����}\�B�g�UG6�E�R?�.mm#ō�҅H��3��݈��b�o�*��x���:�H'��c"�ϋ��>�hNש�iC�HoJ&fJ/�y�~l����I�Ņ�O�&~j���nC��?���HN��J��a��K�ըO�fO�e��r��18��zf���q0\��5�$X+���uq��r�LG�PAC�Ӻ��b�LІe\��(	q���_EV{��@s��Z��Hï�.�������A�k}�I2�	 �KE��4�u�]�%/��Ƿ�p��DJY'8��j>��L��K`Ä
�t�ֹ{[Y-<欚�U�P1t��O��SA�"���dG�B�
}�kuE<��9i�"��a9�'Xj�x��Ԡ	��D�8zx�w=���p_�l��&������den����VH6�t�2'���^L��PtșS���ϓ(�ݙB�	�߆��ÜuMdw�6��N�Kv�"��;奝+Ii�a��\���_���AD�PУ"dqi܈
���?qZ��.U-�u�� 4��;���H��QW3�o��DQA7r �
^��~n�cEPԗ��+A;,��:.?��O�@�-���{g�#��F�/�����e�nf%q�Į�S\wN以��<4���H�)}���=�4NMEM-��{�t��X�8G���¼sY��"�.0���˾���	��(��Y���3AX��d�*)���975���s�u'x�f����z��t�Ca��)�x��c��<�Xߛ����3g!���g��)�69�����B3��2�����&oo�S� AB���qŎ�Գ8K��텣�s'�H`�lc�YK=CV@W-~ҭ�1��:��˓�I!�����M���*����.`�%�ՆF
�z�.�&|̤�/o��+�p�.�"����u��^��͵�jHD8��֕"�}���g��r�[�Y��b���b�7���I�u�="�C�V=�Rϭ�\QRUrE�[?�:�(�� �Ɉ�ȁ}��G���4���I���.�XJ�l���G�����Lu�R�����Џ�M�nq��q��&nI8�e�uj��p�!�=j��ȎX�ze�ѝ��}��-�K �->u�c���$����5cu��轺M�	�!�#��1ibF�T+qA�0e��6���
����@e�I�������K��dO�1�8ek�5g�\�&��ՔXn�,�OXs�ѫpY�)����(&<��h�@�*uOp���>���|��W�tP��Z˸��{\ wmX�hŨn#
X0���j�'�VЖ������������T��Μ�/��I�2�G��^�˕j����:r����@XD��6K��~�.ԋN��j��������=N#"������+V�"od�Fm��yI��kB���2��!|�:����|l��k���@��2�p��Rҁ�=��K��3�m�r7M�X����{�Uj\ozd�z��0�|��F��;7�T��r�'xOy��M���.��xЇ�h�>V�4�nl��jΉƿ��Ƚ��>k�#��Լ��i����~3��T�q��N�h"���OE�#bVn= c�GĖx�,��=!6J-Xz"� 8��L'W���5 ���n���4g^�)чe��/���#���b���~ї�˭w���T(�Xd%�4��5��m�\��>a�F_�y��h�rŲ��;�c����f�țO�V��)P\�[F[[cD�`|���)����]��C6,� m	�8�C'����ϛue�<��4S�^7bW�RPA�z��~p��8�]��K�4��%�EOUw\J�>9��,��#T���n����`��g)��s�N� ��erޡ��*C��N��EP���tw�Xe�R��j�Wʱ��SS��G��0**��2�a��a�(�Z�Z�����Z!hr��u@ϰ�Fço&�0���c`O�١��5�J��@��O��u���:6��+��*D��M{�6��
��⣀ S�� �E���lQm�����2_��P�
I���f�rAR�Q��i���-�=�u�U���.4�h��{�?��[������gvizA��GּY-�K�}�D32�O>Y�y���'�	~#�R�O�cc��.��S�k�����vu ڐ�K�96{M!�	�\.ݯ-m�i�'�-��J[U~�ߞN'Ӿ�5}�p��,on@�K�$�;�l�k��p��3��(�ރ�Ys��u|��d���Vd��#�Z����n$���)���^\d:���(��%U�+�� ܾ)��4<٪�����f�o����tx��1?�S.��`�9���-=���h���-#���c�h�3����K�ba�.�����{l
<E-nN?1K� ��⎪U�U��-�z�
��OB�bT���] Y+O=�j�Vh�>�_�2GL��������!s�޼�mma�R�F%�¯/�@�}�_�%�=Y7�;a�&���P�-E��4F�8��&f���#�H]��v��{G�dK�n��W_
̯��'E�\$9^�<UW�!�lD�6X�fW��Qw�F݅!!��-?��ـFJ�A�^��:j�7�ɘ�X =���:���21S����\4�qw���vÆ�q�%,U��u�*��S9�f�Y��1��產+�q����=d]��v���9�4b]0)�NmH�"
��q���p������P��W�T���˾A��W-�L\����\�W��bJ����;t��D�W@d�x9����U3r�ClM@XF�ѻ9n�	�=c��������考��_:պ�K)#Zp��8��<@�T�*g{���&iN�K\���������l�~�+Y�L%�Ar���4��'��Y��}-�� �@�I�˂�ۣS�/t8=�<*GhT��������jE�h�+>�����K}��5>zx�a>����nӾ��¥Q�f㖶�����<L��z�7���j�z��5���X-�Cb��J�|#�aԥwJm,��sM���m�Ɖ:~n�f��v�Y	� �f��Ç ��Kh3���I��r�nq���'N�p9U�)j�=���<��S����S;0\-��&x���W�V]��+��[W�ē]v�����x�7-��U�{���I$K&�ܥ�=/�\�o�ٙ��
��z�T���G�Ѧ�Vl��	�h藀����y��8�XkA��~�4��_\���w�����D9ci���!�Cӕ^&gY���q�BC��.��r2֌�6�2��� �WXbLš�Q���=�_B&urtIr7c;�\g�귊]�ᙶ�r.)>a��;x��~ɿ�a�� /?��,�h�ݾ�%%D ¯o�jNg�|"�?�DP�tC�uB�#1���Q=�i�p�=��k��0��"T��L��k @o[aтf0�g+؄���p��Q;�ˣ*�]�	,J,�*~9)0.Ȥ����gB��D��+E�D6��5��0��F�[��9:���1:�"��������9���H�G`t�b�\(��:��Tã&���-��������ܶ�s3K*���NB�9�I��գ�&7?����|z�3\X�ǚ�n�j�T��PC���a����)Z��A}��wY�� �h	�:��U��>��,���Ԟ2�u�>��|uH��(6{8$����w�I��Z@D���zw
��Ӭ&���Z�n�"v��JU����A�p>/�!
w,�sA���}���8�$S�����	,������kl�o~D���R���	\펧�<� W>h ���fz��jWPxze3��<����MV�Xkܙ2���7�_	D���6j����!AF��e��,^F�rh#�Ȣ����\����m�=��po����^R�C@E�w��z$��,���L�\ꎍ�M�:(q�����צ�|���`?�_`� eGNV�aE���8�+,^�($��潆֟�%2ziƔ�����jV򴞇��u�UnoE��#�Q�l݃�i���S`�-?>��$׋my��t�)����h.�g���d���46m�R��>ZS�[��8!z���*9�S�]BE��M�r���0k�
j��s9�|�� urw��Q8qB7!�7x�F��K z|�ɮ��b�0�V��-4���rA�
;�p�Z�/}*�q(�Z���5��`֍c����*�?	aU���^��v� ����%��Ʊ��y�?Mn�Cg������93?��9�������t�Y��$��@W���1����	�KN�]�������}��̯����
_B�$G ^��N�����12,�4��j*^�0o����� U���<�BY����$Z�(��S6�60����1,!���`��t���Oe�sE�U1d� �m�e'F9���"�m��R[�/c2�L��L4F\^�u8���TD?�םXjTsk��.ǽ��l�+�
��Nh�r�������O�o-�6��5ſR��ᨫ�x������Qd@])�[�W��A�u��|��!�{���J(����X�f�p��\�mN/���FՉl0�e�ԡ�2Ϛ��d
����M8�8���*��tI}�%��+�Dp`PJ��К�Ɉ��3*[�y(@��{m��I�;(:#�4�W���"��1͟�&�7��n[��}��+��"���͔��!�l�-\C���鴜��S@�P�7�q��p�Ϊ�p�!ǥG��Dk;�L���-ל�=|�����������Q����W/]i�X�}�/k�F(��af~[a�y�D��B��#���i�f貑��@���ݎ�����g�o�3�I�N�����r��@L�N�ԴeK�:��<Bo=�򎳫DNR��z[�'m�#��ҫ{v�G�J�f&Bm�P�c�F��`)dXDb$X(��%'#+��7Չ`!԰�HX.o�����Fq�1�-���J��"Wg�M1o�f�4���|
˲��Q��~���:$;"s�U���J)��k�Ȝ�L�S���އ�I��W]2���3����ίj��e���kk=�ht�S]����@A2�ɅMK����H���s�����X��y*�{���	v�Cv��
�,�A$���/k
����#RY�w�`�6 ��KnA���q�Z���L�o��Q!p�&G���N�փq���Ú-r��ò��8���ڑ�-�k{�4e�������Ŷ���b�z��p@���&���J�}ͨ�@����]��i��<�YW��x,ܺ�z�[��dG�F��,#H9�3�2��j�q� ��	��˺���w�縕
�+��b�B=O�Φw��NU!AO�~"���DF���U_����s�{¸�)�fQ�"I�Q#rٽMWqT���G�t��I���zO�C��